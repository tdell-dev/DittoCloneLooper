module ROM( input [16-1:0] addr, output reg [31:0] outdata );
	always@(*) begin
		case( addr )
			0: outdata = 32'd65536;
			1: outdata = 32'd65535;
			2: outdata = 32'd65534;
			3: outdata = 32'd65533;
			4: outdata = 32'd65532;
			5: outdata = 32'd65531;
			6: outdata = 32'd65530;
			7: outdata = 32'd65529;
			8: outdata = 32'd65528;
			9: outdata = 32'd65527;
			10: outdata = 32'd65526;
			11: outdata = 32'd65525;
			12: outdata = 32'd65524;
			13: outdata = 32'd65523;
			14: outdata = 32'd65522;
			15: outdata = 32'd65521;
			16: outdata = 32'd65520;
			17: outdata = 32'd65519;
			18: outdata = 32'd65518;
			19: outdata = 32'd65517;
			20: outdata = 32'd65516;
			21: outdata = 32'd65515;
			22: outdata = 32'd65514;
			23: outdata = 32'd65513;
			24: outdata = 32'd65512;
			25: outdata = 32'd65511;
			26: outdata = 32'd65510;
			27: outdata = 32'd65509;
			28: outdata = 32'd65508;
			29: outdata = 32'd65507;
			30: outdata = 32'd65506;
			31: outdata = 32'd65505;
			32: outdata = 32'd65504;
			33: outdata = 32'd65503;
			34: outdata = 32'd65502;
			35: outdata = 32'd65501;
			36: outdata = 32'd65500;
			37: outdata = 32'd65499;
			38: outdata = 32'd65498;
			39: outdata = 32'd65497;
			40: outdata = 32'd65496;
			41: outdata = 32'd65495;
			42: outdata = 32'd65494;
			43: outdata = 32'd65493;
			44: outdata = 32'd65492;
			45: outdata = 32'd65491;
			46: outdata = 32'd65490;
			47: outdata = 32'd65489;
			48: outdata = 32'd65488;
			49: outdata = 32'd65487;
			50: outdata = 32'd65486;
			51: outdata = 32'd65485;
			52: outdata = 32'd65484;
			53: outdata = 32'd65483;
			54: outdata = 32'd65482;
			55: outdata = 32'd65481;
			56: outdata = 32'd65480;
			57: outdata = 32'd65479;
			58: outdata = 32'd65478;
			59: outdata = 32'd65477;
			60: outdata = 32'd65476;
			61: outdata = 32'd65475;
			62: outdata = 32'd65474;
			63: outdata = 32'd65473;
			64: outdata = 32'd65472;
			65: outdata = 32'd65471;
			66: outdata = 32'd65470;
			67: outdata = 32'd65469;
			68: outdata = 32'd65468;
			69: outdata = 32'd65467;
			70: outdata = 32'd65466;
			71: outdata = 32'd65465;
			72: outdata = 32'd65464;
			73: outdata = 32'd65463;
			74: outdata = 32'd65462;
			75: outdata = 32'd65461;
			76: outdata = 32'd65460;
			77: outdata = 32'd65459;
			78: outdata = 32'd65458;
			79: outdata = 32'd65457;
			80: outdata = 32'd65456;
			81: outdata = 32'd65455;
			82: outdata = 32'd65454;
			83: outdata = 32'd65453;
			84: outdata = 32'd65452;
			85: outdata = 32'd65451;
			86: outdata = 32'd65450;
			87: outdata = 32'd65449;
			88: outdata = 32'd65448;
			89: outdata = 32'd65447;
			90: outdata = 32'd65446;
			91: outdata = 32'd65445;
			92: outdata = 32'd65444;
			93: outdata = 32'd65443;
			94: outdata = 32'd65442;
			95: outdata = 32'd65441;
			96: outdata = 32'd65440;
			97: outdata = 32'd65439;
			98: outdata = 32'd65438;
			99: outdata = 32'd65437;
			100: outdata = 32'd65436;
			101: outdata = 32'd65435;
			102: outdata = 32'd65434;
			103: outdata = 32'd65433;
			104: outdata = 32'd65432;
			105: outdata = 32'd65431;
			106: outdata = 32'd65430;
			107: outdata = 32'd65429;
			108: outdata = 32'd65428;
			109: outdata = 32'd65427;
			110: outdata = 32'd65426;
			111: outdata = 32'd65425;
			112: outdata = 32'd65424;
			113: outdata = 32'd65423;
			114: outdata = 32'd65422;
			115: outdata = 32'd65421;
			116: outdata = 32'd65420;
			117: outdata = 32'd65419;
			118: outdata = 32'd65418;
			119: outdata = 32'd65417;
			120: outdata = 32'd65416;
			121: outdata = 32'd65415;
			122: outdata = 32'd65414;
			123: outdata = 32'd65413;
			124: outdata = 32'd65412;
			125: outdata = 32'd65411;
			126: outdata = 32'd65410;
			127: outdata = 32'd65409;
			128: outdata = 32'd65408;
			129: outdata = 32'd65407;
			130: outdata = 32'd65406;
			131: outdata = 32'd65405;
			132: outdata = 32'd65404;
			133: outdata = 32'd65403;
			134: outdata = 32'd65402;
			135: outdata = 32'd65401;
			136: outdata = 32'd65400;
			137: outdata = 32'd65399;
			138: outdata = 32'd65398;
			139: outdata = 32'd65397;
			140: outdata = 32'd65396;
			141: outdata = 32'd65395;
			142: outdata = 32'd65394;
			143: outdata = 32'd65393;
			144: outdata = 32'd65392;
			145: outdata = 32'd65391;
			146: outdata = 32'd65390;
			147: outdata = 32'd65389;
			148: outdata = 32'd65388;
			149: outdata = 32'd65387;
			150: outdata = 32'd65386;
			151: outdata = 32'd65385;
			152: outdata = 32'd65384;
			153: outdata = 32'd65383;
			154: outdata = 32'd65382;
			155: outdata = 32'd65381;
			156: outdata = 32'd65380;
			157: outdata = 32'd65379;
			158: outdata = 32'd65378;
			159: outdata = 32'd65377;
			160: outdata = 32'd65376;
			161: outdata = 32'd65375;
			162: outdata = 32'd65374;
			163: outdata = 32'd65373;
			164: outdata = 32'd65372;
			165: outdata = 32'd65371;
			166: outdata = 32'd65370;
			167: outdata = 32'd65369;
			168: outdata = 32'd65368;
			169: outdata = 32'd65367;
			170: outdata = 32'd65366;
			171: outdata = 32'd65365;
			172: outdata = 32'd65364;
			173: outdata = 32'd65363;
			174: outdata = 32'd65362;
			175: outdata = 32'd65361;
			176: outdata = 32'd65360;
			177: outdata = 32'd65359;
			178: outdata = 32'd65358;
			179: outdata = 32'd65357;
			180: outdata = 32'd65356;
			181: outdata = 32'd65355;
			182: outdata = 32'd65354;
			183: outdata = 32'd65353;
			184: outdata = 32'd65352;
			185: outdata = 32'd65351;
			186: outdata = 32'd65350;
			187: outdata = 32'd65349;
			188: outdata = 32'd65348;
			189: outdata = 32'd65347;
			190: outdata = 32'd65346;
			191: outdata = 32'd65345;
			192: outdata = 32'd65344;
			193: outdata = 32'd65343;
			194: outdata = 32'd65342;
			195: outdata = 32'd65341;
			196: outdata = 32'd65340;
			197: outdata = 32'd65339;
			198: outdata = 32'd65338;
			199: outdata = 32'd65337;
			200: outdata = 32'd65336;
			201: outdata = 32'd65335;
			202: outdata = 32'd65334;
			203: outdata = 32'd65333;
			204: outdata = 32'd65332;
			205: outdata = 32'd65331;
			206: outdata = 32'd65330;
			207: outdata = 32'd65329;
			208: outdata = 32'd65328;
			209: outdata = 32'd65327;
			210: outdata = 32'd65326;
			211: outdata = 32'd65325;
			212: outdata = 32'd65324;
			213: outdata = 32'd65323;
			214: outdata = 32'd65322;
			215: outdata = 32'd65321;
			216: outdata = 32'd65320;
			217: outdata = 32'd65319;
			218: outdata = 32'd65318;
			219: outdata = 32'd65317;
			220: outdata = 32'd65316;
			221: outdata = 32'd65315;
			222: outdata = 32'd65314;
			223: outdata = 32'd65313;
			224: outdata = 32'd65312;
			225: outdata = 32'd65311;
			226: outdata = 32'd65310;
			227: outdata = 32'd65309;
			228: outdata = 32'd65308;
			229: outdata = 32'd65307;
			230: outdata = 32'd65306;
			231: outdata = 32'd65305;
			232: outdata = 32'd65304;
			233: outdata = 32'd65303;
			234: outdata = 32'd65302;
			235: outdata = 32'd65301;
			236: outdata = 32'd65300;
			237: outdata = 32'd65299;
			238: outdata = 32'd65298;
			239: outdata = 32'd65297;
			240: outdata = 32'd65296;
			241: outdata = 32'd65295;
			242: outdata = 32'd65294;
			243: outdata = 32'd65293;
			244: outdata = 32'd65292;
			245: outdata = 32'd65291;
			246: outdata = 32'd65290;
			247: outdata = 32'd65289;
			248: outdata = 32'd65288;
			249: outdata = 32'd65287;
			250: outdata = 32'd65286;
			251: outdata = 32'd65285;
			252: outdata = 32'd65284;
			253: outdata = 32'd65283;
			254: outdata = 32'd65282;
			255: outdata = 32'd65281;
			256: outdata = 32'd65280;
			257: outdata = 32'd65279;
			258: outdata = 32'd65278;
			259: outdata = 32'd65277;
			260: outdata = 32'd65276;
			261: outdata = 32'd65275;
			262: outdata = 32'd65274;
			263: outdata = 32'd65273;
			264: outdata = 32'd65272;
			265: outdata = 32'd65271;
			266: outdata = 32'd65270;
			267: outdata = 32'd65269;
			268: outdata = 32'd65268;
			269: outdata = 32'd65267;
			270: outdata = 32'd65266;
			271: outdata = 32'd65265;
			272: outdata = 32'd65264;
			273: outdata = 32'd65263;
			274: outdata = 32'd65262;
			275: outdata = 32'd65261;
			276: outdata = 32'd65260;
			277: outdata = 32'd65259;
			278: outdata = 32'd65258;
			279: outdata = 32'd65257;
			280: outdata = 32'd65256;
			281: outdata = 32'd65255;
			282: outdata = 32'd65254;
			283: outdata = 32'd65253;
			284: outdata = 32'd65252;
			285: outdata = 32'd65251;
			286: outdata = 32'd65250;
			287: outdata = 32'd65249;
			288: outdata = 32'd65248;
			289: outdata = 32'd65247;
			290: outdata = 32'd65246;
			291: outdata = 32'd65245;
			292: outdata = 32'd65244;
			293: outdata = 32'd65243;
			294: outdata = 32'd65242;
			295: outdata = 32'd65241;
			296: outdata = 32'd65240;
			297: outdata = 32'd65239;
			298: outdata = 32'd65238;
			299: outdata = 32'd65237;
			300: outdata = 32'd65236;
			301: outdata = 32'd65235;
			302: outdata = 32'd65234;
			303: outdata = 32'd65233;
			304: outdata = 32'd65232;
			305: outdata = 32'd65231;
			306: outdata = 32'd65230;
			307: outdata = 32'd65229;
			308: outdata = 32'd65228;
			309: outdata = 32'd65227;
			310: outdata = 32'd65226;
			311: outdata = 32'd65225;
			312: outdata = 32'd65224;
			313: outdata = 32'd65223;
			314: outdata = 32'd65222;
			315: outdata = 32'd65221;
			316: outdata = 32'd65220;
			317: outdata = 32'd65219;
			318: outdata = 32'd65218;
			319: outdata = 32'd65217;
			320: outdata = 32'd65216;
			321: outdata = 32'd65215;
			322: outdata = 32'd65214;
			323: outdata = 32'd65213;
			324: outdata = 32'd65212;
			325: outdata = 32'd65211;
			326: outdata = 32'd65210;
			327: outdata = 32'd65209;
			328: outdata = 32'd65208;
			329: outdata = 32'd65207;
			330: outdata = 32'd65206;
			331: outdata = 32'd65205;
			332: outdata = 32'd65204;
			333: outdata = 32'd65203;
			334: outdata = 32'd65202;
			335: outdata = 32'd65201;
			336: outdata = 32'd65200;
			337: outdata = 32'd65199;
			338: outdata = 32'd65198;
			339: outdata = 32'd65197;
			340: outdata = 32'd65196;
			341: outdata = 32'd65195;
			342: outdata = 32'd65194;
			343: outdata = 32'd65193;
			344: outdata = 32'd65192;
			345: outdata = 32'd65191;
			346: outdata = 32'd65190;
			347: outdata = 32'd65189;
			348: outdata = 32'd65188;
			349: outdata = 32'd65187;
			350: outdata = 32'd65186;
			351: outdata = 32'd65185;
			352: outdata = 32'd65184;
			353: outdata = 32'd65183;
			354: outdata = 32'd65182;
			355: outdata = 32'd65181;
			356: outdata = 32'd65180;
			357: outdata = 32'd65179;
			358: outdata = 32'd65178;
			359: outdata = 32'd65177;
			360: outdata = 32'd65176;
			361: outdata = 32'd65175;
			362: outdata = 32'd65174;
			363: outdata = 32'd65173;
			364: outdata = 32'd65172;
			365: outdata = 32'd65171;
			366: outdata = 32'd65170;
			367: outdata = 32'd65169;
			368: outdata = 32'd65168;
			369: outdata = 32'd65167;
			370: outdata = 32'd65166;
			371: outdata = 32'd65165;
			372: outdata = 32'd65164;
			373: outdata = 32'd65163;
			374: outdata = 32'd65162;
			375: outdata = 32'd65161;
			376: outdata = 32'd65160;
			377: outdata = 32'd65159;
			378: outdata = 32'd65158;
			379: outdata = 32'd65157;
			380: outdata = 32'd65156;
			381: outdata = 32'd65155;
			382: outdata = 32'd65154;
			383: outdata = 32'd65153;
			384: outdata = 32'd65152;
			385: outdata = 32'd65151;
			386: outdata = 32'd65150;
			387: outdata = 32'd65149;
			388: outdata = 32'd65148;
			389: outdata = 32'd65147;
			390: outdata = 32'd65146;
			391: outdata = 32'd65145;
			392: outdata = 32'd65144;
			393: outdata = 32'd65143;
			394: outdata = 32'd65142;
			395: outdata = 32'd65141;
			396: outdata = 32'd65140;
			397: outdata = 32'd65139;
			398: outdata = 32'd65138;
			399: outdata = 32'd65137;
			400: outdata = 32'd65136;
			401: outdata = 32'd65135;
			402: outdata = 32'd65134;
			403: outdata = 32'd65133;
			404: outdata = 32'd65132;
			405: outdata = 32'd65131;
			406: outdata = 32'd65130;
			407: outdata = 32'd65129;
			408: outdata = 32'd65128;
			409: outdata = 32'd65127;
			410: outdata = 32'd65126;
			411: outdata = 32'd65125;
			412: outdata = 32'd65124;
			413: outdata = 32'd65123;
			414: outdata = 32'd65122;
			415: outdata = 32'd65121;
			416: outdata = 32'd65120;
			417: outdata = 32'd65119;
			418: outdata = 32'd65118;
			419: outdata = 32'd65117;
			420: outdata = 32'd65116;
			421: outdata = 32'd65115;
			422: outdata = 32'd65114;
			423: outdata = 32'd65113;
			424: outdata = 32'd65112;
			425: outdata = 32'd65111;
			426: outdata = 32'd65110;
			427: outdata = 32'd65109;
			428: outdata = 32'd65108;
			429: outdata = 32'd65107;
			430: outdata = 32'd65106;
			431: outdata = 32'd65105;
			432: outdata = 32'd65104;
			433: outdata = 32'd65103;
			434: outdata = 32'd65102;
			435: outdata = 32'd65101;
			436: outdata = 32'd65100;
			437: outdata = 32'd65099;
			438: outdata = 32'd65098;
			439: outdata = 32'd65097;
			440: outdata = 32'd65096;
			441: outdata = 32'd65095;
			442: outdata = 32'd65094;
			443: outdata = 32'd65093;
			444: outdata = 32'd65092;
			445: outdata = 32'd65091;
			446: outdata = 32'd65090;
			447: outdata = 32'd65089;
			448: outdata = 32'd65088;
			449: outdata = 32'd65087;
			450: outdata = 32'd65086;
			451: outdata = 32'd65085;
			452: outdata = 32'd65084;
			453: outdata = 32'd65083;
			454: outdata = 32'd65082;
			455: outdata = 32'd65081;
			456: outdata = 32'd65080;
			457: outdata = 32'd65079;
			458: outdata = 32'd65078;
			459: outdata = 32'd65077;
			460: outdata = 32'd65076;
			461: outdata = 32'd65075;
			462: outdata = 32'd65074;
			463: outdata = 32'd65073;
			464: outdata = 32'd65072;
			465: outdata = 32'd65071;
			466: outdata = 32'd65070;
			467: outdata = 32'd65069;
			468: outdata = 32'd65068;
			469: outdata = 32'd65067;
			470: outdata = 32'd65066;
			471: outdata = 32'd65065;
			472: outdata = 32'd65064;
			473: outdata = 32'd65063;
			474: outdata = 32'd65062;
			475: outdata = 32'd65061;
			476: outdata = 32'd65060;
			477: outdata = 32'd65059;
			478: outdata = 32'd65058;
			479: outdata = 32'd65057;
			480: outdata = 32'd65056;
			481: outdata = 32'd65055;
			482: outdata = 32'd65054;
			483: outdata = 32'd65053;
			484: outdata = 32'd65052;
			485: outdata = 32'd65051;
			486: outdata = 32'd65050;
			487: outdata = 32'd65049;
			488: outdata = 32'd65048;
			489: outdata = 32'd65047;
			490: outdata = 32'd65046;
			491: outdata = 32'd65045;
			492: outdata = 32'd65044;
			493: outdata = 32'd65043;
			494: outdata = 32'd65042;
			495: outdata = 32'd65041;
			496: outdata = 32'd65040;
			497: outdata = 32'd65039;
			498: outdata = 32'd65038;
			499: outdata = 32'd65037;
			500: outdata = 32'd65036;
			501: outdata = 32'd65035;
			502: outdata = 32'd65034;
			503: outdata = 32'd65033;
			504: outdata = 32'd65032;
			505: outdata = 32'd65031;
			506: outdata = 32'd65030;
			507: outdata = 32'd65029;
			508: outdata = 32'd65028;
			509: outdata = 32'd65027;
			510: outdata = 32'd65026;
			511: outdata = 32'd65025;
			512: outdata = 32'd65024;
			513: outdata = 32'd65023;
			514: outdata = 32'd65022;
			515: outdata = 32'd65021;
			516: outdata = 32'd65020;
			517: outdata = 32'd65019;
			518: outdata = 32'd65018;
			519: outdata = 32'd65017;
			520: outdata = 32'd65016;
			521: outdata = 32'd65015;
			522: outdata = 32'd65014;
			523: outdata = 32'd65013;
			524: outdata = 32'd65012;
			525: outdata = 32'd65011;
			526: outdata = 32'd65010;
			527: outdata = 32'd65009;
			528: outdata = 32'd65008;
			529: outdata = 32'd65007;
			530: outdata = 32'd65006;
			531: outdata = 32'd65005;
			532: outdata = 32'd65004;
			533: outdata = 32'd65003;
			534: outdata = 32'd65002;
			535: outdata = 32'd65001;
			536: outdata = 32'd65000;
			537: outdata = 32'd64999;
			538: outdata = 32'd64998;
			539: outdata = 32'd64997;
			540: outdata = 32'd64996;
			541: outdata = 32'd64995;
			542: outdata = 32'd64994;
			543: outdata = 32'd64993;
			544: outdata = 32'd64992;
			545: outdata = 32'd64991;
			546: outdata = 32'd64990;
			547: outdata = 32'd64989;
			548: outdata = 32'd64988;
			549: outdata = 32'd64987;
			550: outdata = 32'd64986;
			551: outdata = 32'd64985;
			552: outdata = 32'd64984;
			553: outdata = 32'd64983;
			554: outdata = 32'd64982;
			555: outdata = 32'd64981;
			556: outdata = 32'd64980;
			557: outdata = 32'd64979;
			558: outdata = 32'd64978;
			559: outdata = 32'd64977;
			560: outdata = 32'd64976;
			561: outdata = 32'd64975;
			562: outdata = 32'd64974;
			563: outdata = 32'd64973;
			564: outdata = 32'd64972;
			565: outdata = 32'd64971;
			566: outdata = 32'd64970;
			567: outdata = 32'd64969;
			568: outdata = 32'd64968;
			569: outdata = 32'd64967;
			570: outdata = 32'd64966;
			571: outdata = 32'd64965;
			572: outdata = 32'd64964;
			573: outdata = 32'd64963;
			574: outdata = 32'd64962;
			575: outdata = 32'd64961;
			576: outdata = 32'd64960;
			577: outdata = 32'd64959;
			578: outdata = 32'd64958;
			579: outdata = 32'd64957;
			580: outdata = 32'd64956;
			581: outdata = 32'd64955;
			582: outdata = 32'd64954;
			583: outdata = 32'd64953;
			584: outdata = 32'd64952;
			585: outdata = 32'd64951;
			586: outdata = 32'd64950;
			587: outdata = 32'd64949;
			588: outdata = 32'd64948;
			589: outdata = 32'd64947;
			590: outdata = 32'd64946;
			591: outdata = 32'd64945;
			592: outdata = 32'd64944;
			593: outdata = 32'd64943;
			594: outdata = 32'd64942;
			595: outdata = 32'd64941;
			596: outdata = 32'd64940;
			597: outdata = 32'd64939;
			598: outdata = 32'd64938;
			599: outdata = 32'd64937;
			600: outdata = 32'd64936;
			601: outdata = 32'd64935;
			602: outdata = 32'd64934;
			603: outdata = 32'd64933;
			604: outdata = 32'd64932;
			605: outdata = 32'd64931;
			606: outdata = 32'd64930;
			607: outdata = 32'd64929;
			608: outdata = 32'd64928;
			609: outdata = 32'd64927;
			610: outdata = 32'd64926;
			611: outdata = 32'd64925;
			612: outdata = 32'd64924;
			613: outdata = 32'd64923;
			614: outdata = 32'd64922;
			615: outdata = 32'd64921;
			616: outdata = 32'd64920;
			617: outdata = 32'd64919;
			618: outdata = 32'd64918;
			619: outdata = 32'd64917;
			620: outdata = 32'd64916;
			621: outdata = 32'd64915;
			622: outdata = 32'd64914;
			623: outdata = 32'd64913;
			624: outdata = 32'd64912;
			625: outdata = 32'd64911;
			626: outdata = 32'd64910;
			627: outdata = 32'd64909;
			628: outdata = 32'd64908;
			629: outdata = 32'd64907;
			630: outdata = 32'd64906;
			631: outdata = 32'd64905;
			632: outdata = 32'd64904;
			633: outdata = 32'd64903;
			634: outdata = 32'd64902;
			635: outdata = 32'd64901;
			636: outdata = 32'd64900;
			637: outdata = 32'd64899;
			638: outdata = 32'd64898;
			639: outdata = 32'd64897;
			640: outdata = 32'd64896;
			641: outdata = 32'd64895;
			642: outdata = 32'd64894;
			643: outdata = 32'd64893;
			644: outdata = 32'd64892;
			645: outdata = 32'd64891;
			646: outdata = 32'd64890;
			647: outdata = 32'd64889;
			648: outdata = 32'd64888;
			649: outdata = 32'd64887;
			650: outdata = 32'd64886;
			651: outdata = 32'd64885;
			652: outdata = 32'd64884;
			653: outdata = 32'd64883;
			654: outdata = 32'd64882;
			655: outdata = 32'd64881;
			656: outdata = 32'd64880;
			657: outdata = 32'd64879;
			658: outdata = 32'd64878;
			659: outdata = 32'd64877;
			660: outdata = 32'd64876;
			661: outdata = 32'd64875;
			662: outdata = 32'd64874;
			663: outdata = 32'd64873;
			664: outdata = 32'd64872;
			665: outdata = 32'd64871;
			666: outdata = 32'd64870;
			667: outdata = 32'd64869;
			668: outdata = 32'd64868;
			669: outdata = 32'd64867;
			670: outdata = 32'd64866;
			671: outdata = 32'd64865;
			672: outdata = 32'd64864;
			673: outdata = 32'd64863;
			674: outdata = 32'd64862;
			675: outdata = 32'd64861;
			676: outdata = 32'd64860;
			677: outdata = 32'd64859;
			678: outdata = 32'd64858;
			679: outdata = 32'd64857;
			680: outdata = 32'd64856;
			681: outdata = 32'd64855;
			682: outdata = 32'd64854;
			683: outdata = 32'd64853;
			684: outdata = 32'd64852;
			685: outdata = 32'd64851;
			686: outdata = 32'd64850;
			687: outdata = 32'd64849;
			688: outdata = 32'd64848;
			689: outdata = 32'd64847;
			690: outdata = 32'd64846;
			691: outdata = 32'd64845;
			692: outdata = 32'd64844;
			693: outdata = 32'd64843;
			694: outdata = 32'd64842;
			695: outdata = 32'd64841;
			696: outdata = 32'd64840;
			697: outdata = 32'd64839;
			698: outdata = 32'd64838;
			699: outdata = 32'd64837;
			700: outdata = 32'd64836;
			701: outdata = 32'd64835;
			702: outdata = 32'd64834;
			703: outdata = 32'd64833;
			704: outdata = 32'd64832;
			705: outdata = 32'd64831;
			706: outdata = 32'd64830;
			707: outdata = 32'd64829;
			708: outdata = 32'd64828;
			709: outdata = 32'd64827;
			710: outdata = 32'd64826;
			711: outdata = 32'd64825;
			712: outdata = 32'd64824;
			713: outdata = 32'd64823;
			714: outdata = 32'd64822;
			715: outdata = 32'd64821;
			716: outdata = 32'd64820;
			717: outdata = 32'd64819;
			718: outdata = 32'd64818;
			719: outdata = 32'd64817;
			720: outdata = 32'd64816;
			721: outdata = 32'd64815;
			722: outdata = 32'd64814;
			723: outdata = 32'd64813;
			724: outdata = 32'd64812;
			725: outdata = 32'd64811;
			726: outdata = 32'd64810;
			727: outdata = 32'd64809;
			728: outdata = 32'd64808;
			729: outdata = 32'd64807;
			730: outdata = 32'd64806;
			731: outdata = 32'd64805;
			732: outdata = 32'd64804;
			733: outdata = 32'd64803;
			734: outdata = 32'd64802;
			735: outdata = 32'd64801;
			736: outdata = 32'd64800;
			737: outdata = 32'd64799;
			738: outdata = 32'd64798;
			739: outdata = 32'd64797;
			740: outdata = 32'd64796;
			741: outdata = 32'd64795;
			742: outdata = 32'd64794;
			743: outdata = 32'd64793;
			744: outdata = 32'd64792;
			745: outdata = 32'd64791;
			746: outdata = 32'd64790;
			747: outdata = 32'd64789;
			748: outdata = 32'd64788;
			749: outdata = 32'd64787;
			750: outdata = 32'd64786;
			751: outdata = 32'd64785;
			752: outdata = 32'd64784;
			753: outdata = 32'd64783;
			754: outdata = 32'd64782;
			755: outdata = 32'd64781;
			756: outdata = 32'd64780;
			757: outdata = 32'd64779;
			758: outdata = 32'd64778;
			759: outdata = 32'd64777;
			760: outdata = 32'd64776;
			761: outdata = 32'd64775;
			762: outdata = 32'd64774;
			763: outdata = 32'd64773;
			764: outdata = 32'd64772;
			765: outdata = 32'd64771;
			766: outdata = 32'd64770;
			767: outdata = 32'd64769;
			768: outdata = 32'd64768;
			769: outdata = 32'd64767;
			770: outdata = 32'd64766;
			771: outdata = 32'd64765;
			772: outdata = 32'd64764;
			773: outdata = 32'd64763;
			774: outdata = 32'd64762;
			775: outdata = 32'd64761;
			776: outdata = 32'd64760;
			777: outdata = 32'd64759;
			778: outdata = 32'd64758;
			779: outdata = 32'd64757;
			780: outdata = 32'd64756;
			781: outdata = 32'd64755;
			782: outdata = 32'd64754;
			783: outdata = 32'd64753;
			784: outdata = 32'd64752;
			785: outdata = 32'd64751;
			786: outdata = 32'd64750;
			787: outdata = 32'd64749;
			788: outdata = 32'd64748;
			789: outdata = 32'd64747;
			790: outdata = 32'd64746;
			791: outdata = 32'd64745;
			792: outdata = 32'd64744;
			793: outdata = 32'd64743;
			794: outdata = 32'd64742;
			795: outdata = 32'd64741;
			796: outdata = 32'd64740;
			797: outdata = 32'd64739;
			798: outdata = 32'd64738;
			799: outdata = 32'd64737;
			800: outdata = 32'd64736;
			801: outdata = 32'd64735;
			802: outdata = 32'd64734;
			803: outdata = 32'd64733;
			804: outdata = 32'd64732;
			805: outdata = 32'd64731;
			806: outdata = 32'd64730;
			807: outdata = 32'd64729;
			808: outdata = 32'd64728;
			809: outdata = 32'd64727;
			810: outdata = 32'd64726;
			811: outdata = 32'd64725;
			812: outdata = 32'd64724;
			813: outdata = 32'd64723;
			814: outdata = 32'd64722;
			815: outdata = 32'd64721;
			816: outdata = 32'd64720;
			817: outdata = 32'd64719;
			818: outdata = 32'd64718;
			819: outdata = 32'd64717;
			820: outdata = 32'd64716;
			821: outdata = 32'd64715;
			822: outdata = 32'd64714;
			823: outdata = 32'd64713;
			824: outdata = 32'd64712;
			825: outdata = 32'd64711;
			826: outdata = 32'd64710;
			827: outdata = 32'd64709;
			828: outdata = 32'd64708;
			829: outdata = 32'd64707;
			830: outdata = 32'd64706;
			831: outdata = 32'd64705;
			832: outdata = 32'd64704;
			833: outdata = 32'd64703;
			834: outdata = 32'd64702;
			835: outdata = 32'd64701;
			836: outdata = 32'd64700;
			837: outdata = 32'd64699;
			838: outdata = 32'd64698;
			839: outdata = 32'd64697;
			840: outdata = 32'd64696;
			841: outdata = 32'd64695;
			842: outdata = 32'd64694;
			843: outdata = 32'd64693;
			844: outdata = 32'd64692;
			845: outdata = 32'd64691;
			846: outdata = 32'd64690;
			847: outdata = 32'd64689;
			848: outdata = 32'd64688;
			849: outdata = 32'd64687;
			850: outdata = 32'd64686;
			851: outdata = 32'd64685;
			852: outdata = 32'd64684;
			853: outdata = 32'd64683;
			854: outdata = 32'd64682;
			855: outdata = 32'd64681;
			856: outdata = 32'd64680;
			857: outdata = 32'd64679;
			858: outdata = 32'd64678;
			859: outdata = 32'd64677;
			860: outdata = 32'd64676;
			861: outdata = 32'd64675;
			862: outdata = 32'd64674;
			863: outdata = 32'd64673;
			864: outdata = 32'd64672;
			865: outdata = 32'd64671;
			866: outdata = 32'd64670;
			867: outdata = 32'd64669;
			868: outdata = 32'd64668;
			869: outdata = 32'd64667;
			870: outdata = 32'd64666;
			871: outdata = 32'd64665;
			872: outdata = 32'd64664;
			873: outdata = 32'd64663;
			874: outdata = 32'd64662;
			875: outdata = 32'd64661;
			876: outdata = 32'd64660;
			877: outdata = 32'd64659;
			878: outdata = 32'd64658;
			879: outdata = 32'd64657;
			880: outdata = 32'd64656;
			881: outdata = 32'd64655;
			882: outdata = 32'd64654;
			883: outdata = 32'd64653;
			884: outdata = 32'd64652;
			885: outdata = 32'd64651;
			886: outdata = 32'd64650;
			887: outdata = 32'd64649;
			888: outdata = 32'd64648;
			889: outdata = 32'd64647;
			890: outdata = 32'd64646;
			891: outdata = 32'd64645;
			892: outdata = 32'd64644;
			893: outdata = 32'd64643;
			894: outdata = 32'd64642;
			895: outdata = 32'd64641;
			896: outdata = 32'd64640;
			897: outdata = 32'd64639;
			898: outdata = 32'd64638;
			899: outdata = 32'd64637;
			900: outdata = 32'd64636;
			901: outdata = 32'd64635;
			902: outdata = 32'd64634;
			903: outdata = 32'd64633;
			904: outdata = 32'd64632;
			905: outdata = 32'd64631;
			906: outdata = 32'd64630;
			907: outdata = 32'd64629;
			908: outdata = 32'd64628;
			909: outdata = 32'd64627;
			910: outdata = 32'd64626;
			911: outdata = 32'd64625;
			912: outdata = 32'd64624;
			913: outdata = 32'd64623;
			914: outdata = 32'd64622;
			915: outdata = 32'd64621;
			916: outdata = 32'd64620;
			917: outdata = 32'd64619;
			918: outdata = 32'd64618;
			919: outdata = 32'd64617;
			920: outdata = 32'd64616;
			921: outdata = 32'd64615;
			922: outdata = 32'd64614;
			923: outdata = 32'd64613;
			924: outdata = 32'd64612;
			925: outdata = 32'd64611;
			926: outdata = 32'd64610;
			927: outdata = 32'd64609;
			928: outdata = 32'd64608;
			929: outdata = 32'd64607;
			930: outdata = 32'd64606;
			931: outdata = 32'd64605;
			932: outdata = 32'd64604;
			933: outdata = 32'd64603;
			934: outdata = 32'd64602;
			935: outdata = 32'd64601;
			936: outdata = 32'd64600;
			937: outdata = 32'd64599;
			938: outdata = 32'd64598;
			939: outdata = 32'd64597;
			940: outdata = 32'd64596;
			941: outdata = 32'd64595;
			942: outdata = 32'd64594;
			943: outdata = 32'd64593;
			944: outdata = 32'd64592;
			945: outdata = 32'd64591;
			946: outdata = 32'd64590;
			947: outdata = 32'd64589;
			948: outdata = 32'd64588;
			949: outdata = 32'd64587;
			950: outdata = 32'd64586;
			951: outdata = 32'd64585;
			952: outdata = 32'd64584;
			953: outdata = 32'd64583;
			954: outdata = 32'd64582;
			955: outdata = 32'd64581;
			956: outdata = 32'd64580;
			957: outdata = 32'd64579;
			958: outdata = 32'd64578;
			959: outdata = 32'd64577;
			960: outdata = 32'd64576;
			961: outdata = 32'd64575;
			962: outdata = 32'd64574;
			963: outdata = 32'd64573;
			964: outdata = 32'd64572;
			965: outdata = 32'd64571;
			966: outdata = 32'd64570;
			967: outdata = 32'd64569;
			968: outdata = 32'd64568;
			969: outdata = 32'd64567;
			970: outdata = 32'd64566;
			971: outdata = 32'd64565;
			972: outdata = 32'd64564;
			973: outdata = 32'd64563;
			974: outdata = 32'd64562;
			975: outdata = 32'd64561;
			976: outdata = 32'd64560;
			977: outdata = 32'd64559;
			978: outdata = 32'd64558;
			979: outdata = 32'd64557;
			980: outdata = 32'd64556;
			981: outdata = 32'd64555;
			982: outdata = 32'd64554;
			983: outdata = 32'd64553;
			984: outdata = 32'd64552;
			985: outdata = 32'd64551;
			986: outdata = 32'd64550;
			987: outdata = 32'd64549;
			988: outdata = 32'd64548;
			989: outdata = 32'd64547;
			990: outdata = 32'd64546;
			991: outdata = 32'd64545;
			992: outdata = 32'd64544;
			993: outdata = 32'd64543;
			994: outdata = 32'd64542;
			995: outdata = 32'd64541;
			996: outdata = 32'd64540;
			997: outdata = 32'd64539;
			998: outdata = 32'd64538;
			999: outdata = 32'd64537;
			1000: outdata = 32'd64536;
			1001: outdata = 32'd64535;
			1002: outdata = 32'd64534;
			1003: outdata = 32'd64533;
			1004: outdata = 32'd64532;
			1005: outdata = 32'd64531;
			1006: outdata = 32'd64530;
			1007: outdata = 32'd64529;
			1008: outdata = 32'd64528;
			1009: outdata = 32'd64527;
			1010: outdata = 32'd64526;
			1011: outdata = 32'd64525;
			1012: outdata = 32'd64524;
			1013: outdata = 32'd64523;
			1014: outdata = 32'd64522;
			1015: outdata = 32'd64521;
			1016: outdata = 32'd64520;
			1017: outdata = 32'd64519;
			1018: outdata = 32'd64518;
			1019: outdata = 32'd64517;
			1020: outdata = 32'd64516;
			1021: outdata = 32'd64515;
			1022: outdata = 32'd64514;
			1023: outdata = 32'd64513;
			1024: outdata = 32'd64512;
			1025: outdata = 32'd64511;
			1026: outdata = 32'd64510;
			1027: outdata = 32'd64509;
			1028: outdata = 32'd64508;
			1029: outdata = 32'd64507;
			1030: outdata = 32'd64506;
			1031: outdata = 32'd64505;
			1032: outdata = 32'd64504;
			1033: outdata = 32'd64503;
			1034: outdata = 32'd64502;
			1035: outdata = 32'd64501;
			1036: outdata = 32'd64500;
			1037: outdata = 32'd64499;
			1038: outdata = 32'd64498;
			1039: outdata = 32'd64497;
			1040: outdata = 32'd64496;
			1041: outdata = 32'd64495;
			1042: outdata = 32'd64494;
			1043: outdata = 32'd64493;
			1044: outdata = 32'd64492;
			1045: outdata = 32'd64491;
			1046: outdata = 32'd64490;
			1047: outdata = 32'd64489;
			1048: outdata = 32'd64488;
			1049: outdata = 32'd64487;
			1050: outdata = 32'd64486;
			1051: outdata = 32'd64485;
			1052: outdata = 32'd64484;
			1053: outdata = 32'd64483;
			1054: outdata = 32'd64482;
			1055: outdata = 32'd64481;
			1056: outdata = 32'd64480;
			1057: outdata = 32'd64479;
			1058: outdata = 32'd64478;
			1059: outdata = 32'd64477;
			1060: outdata = 32'd64476;
			1061: outdata = 32'd64475;
			1062: outdata = 32'd64474;
			1063: outdata = 32'd64473;
			1064: outdata = 32'd64472;
			1065: outdata = 32'd64471;
			1066: outdata = 32'd64470;
			1067: outdata = 32'd64469;
			1068: outdata = 32'd64468;
			1069: outdata = 32'd64467;
			1070: outdata = 32'd64466;
			1071: outdata = 32'd64465;
			1072: outdata = 32'd64464;
			1073: outdata = 32'd64463;
			1074: outdata = 32'd64462;
			1075: outdata = 32'd64461;
			1076: outdata = 32'd64460;
			1077: outdata = 32'd64459;
			1078: outdata = 32'd64458;
			1079: outdata = 32'd64457;
			1080: outdata = 32'd64456;
			1081: outdata = 32'd64455;
			1082: outdata = 32'd64454;
			1083: outdata = 32'd64453;
			1084: outdata = 32'd64452;
			1085: outdata = 32'd64451;
			1086: outdata = 32'd64450;
			1087: outdata = 32'd64449;
			1088: outdata = 32'd64448;
			1089: outdata = 32'd64447;
			1090: outdata = 32'd64446;
			1091: outdata = 32'd64445;
			1092: outdata = 32'd64444;
			1093: outdata = 32'd64443;
			1094: outdata = 32'd64442;
			1095: outdata = 32'd64441;
			1096: outdata = 32'd64440;
			1097: outdata = 32'd64439;
			1098: outdata = 32'd64438;
			1099: outdata = 32'd64437;
			1100: outdata = 32'd64436;
			1101: outdata = 32'd64435;
			1102: outdata = 32'd64434;
			1103: outdata = 32'd64433;
			1104: outdata = 32'd64432;
			1105: outdata = 32'd64431;
			1106: outdata = 32'd64430;
			1107: outdata = 32'd64429;
			1108: outdata = 32'd64428;
			1109: outdata = 32'd64427;
			1110: outdata = 32'd64426;
			1111: outdata = 32'd64425;
			1112: outdata = 32'd64424;
			1113: outdata = 32'd64423;
			1114: outdata = 32'd64422;
			1115: outdata = 32'd64421;
			1116: outdata = 32'd64420;
			1117: outdata = 32'd64419;
			1118: outdata = 32'd64418;
			1119: outdata = 32'd64417;
			1120: outdata = 32'd64416;
			1121: outdata = 32'd64415;
			1122: outdata = 32'd64414;
			1123: outdata = 32'd64413;
			1124: outdata = 32'd64412;
			1125: outdata = 32'd64411;
			1126: outdata = 32'd64410;
			1127: outdata = 32'd64409;
			1128: outdata = 32'd64408;
			1129: outdata = 32'd64407;
			1130: outdata = 32'd64406;
			1131: outdata = 32'd64405;
			1132: outdata = 32'd64404;
			1133: outdata = 32'd64403;
			1134: outdata = 32'd64402;
			1135: outdata = 32'd64401;
			1136: outdata = 32'd64400;
			1137: outdata = 32'd64399;
			1138: outdata = 32'd64398;
			1139: outdata = 32'd64397;
			1140: outdata = 32'd64396;
			1141: outdata = 32'd64395;
			1142: outdata = 32'd64394;
			1143: outdata = 32'd64393;
			1144: outdata = 32'd64392;
			1145: outdata = 32'd64391;
			1146: outdata = 32'd64390;
			1147: outdata = 32'd64389;
			1148: outdata = 32'd64388;
			1149: outdata = 32'd64387;
			1150: outdata = 32'd64386;
			1151: outdata = 32'd64385;
			1152: outdata = 32'd64384;
			1153: outdata = 32'd64383;
			1154: outdata = 32'd64382;
			1155: outdata = 32'd64381;
			1156: outdata = 32'd64380;
			1157: outdata = 32'd64379;
			1158: outdata = 32'd64378;
			1159: outdata = 32'd64377;
			1160: outdata = 32'd64376;
			1161: outdata = 32'd64375;
			1162: outdata = 32'd64374;
			1163: outdata = 32'd64373;
			1164: outdata = 32'd64372;
			1165: outdata = 32'd64371;
			1166: outdata = 32'd64370;
			1167: outdata = 32'd64369;
			1168: outdata = 32'd64368;
			1169: outdata = 32'd64367;
			1170: outdata = 32'd64366;
			1171: outdata = 32'd64365;
			1172: outdata = 32'd64364;
			1173: outdata = 32'd64363;
			1174: outdata = 32'd64362;
			1175: outdata = 32'd64361;
			1176: outdata = 32'd64360;
			1177: outdata = 32'd64359;
			1178: outdata = 32'd64358;
			1179: outdata = 32'd64357;
			1180: outdata = 32'd64356;
			1181: outdata = 32'd64355;
			1182: outdata = 32'd64354;
			1183: outdata = 32'd64353;
			1184: outdata = 32'd64352;
			1185: outdata = 32'd64351;
			1186: outdata = 32'd64350;
			1187: outdata = 32'd64349;
			1188: outdata = 32'd64348;
			1189: outdata = 32'd64347;
			1190: outdata = 32'd64346;
			1191: outdata = 32'd64345;
			1192: outdata = 32'd64344;
			1193: outdata = 32'd64343;
			1194: outdata = 32'd64342;
			1195: outdata = 32'd64341;
			1196: outdata = 32'd64340;
			1197: outdata = 32'd64339;
			1198: outdata = 32'd64338;
			1199: outdata = 32'd64337;
			1200: outdata = 32'd64336;
			1201: outdata = 32'd64335;
			1202: outdata = 32'd64334;
			1203: outdata = 32'd64333;
			1204: outdata = 32'd64332;
			1205: outdata = 32'd64331;
			1206: outdata = 32'd64330;
			1207: outdata = 32'd64329;
			1208: outdata = 32'd64328;
			1209: outdata = 32'd64327;
			1210: outdata = 32'd64326;
			1211: outdata = 32'd64325;
			1212: outdata = 32'd64324;
			1213: outdata = 32'd64323;
			1214: outdata = 32'd64322;
			1215: outdata = 32'd64321;
			1216: outdata = 32'd64320;
			1217: outdata = 32'd64319;
			1218: outdata = 32'd64318;
			1219: outdata = 32'd64317;
			1220: outdata = 32'd64316;
			1221: outdata = 32'd64315;
			1222: outdata = 32'd64314;
			1223: outdata = 32'd64313;
			1224: outdata = 32'd64312;
			1225: outdata = 32'd64311;
			1226: outdata = 32'd64310;
			1227: outdata = 32'd64309;
			1228: outdata = 32'd64308;
			1229: outdata = 32'd64307;
			1230: outdata = 32'd64306;
			1231: outdata = 32'd64305;
			1232: outdata = 32'd64304;
			1233: outdata = 32'd64303;
			1234: outdata = 32'd64302;
			1235: outdata = 32'd64301;
			1236: outdata = 32'd64300;
			1237: outdata = 32'd64299;
			1238: outdata = 32'd64298;
			1239: outdata = 32'd64297;
			1240: outdata = 32'd64296;
			1241: outdata = 32'd64295;
			1242: outdata = 32'd64294;
			1243: outdata = 32'd64293;
			1244: outdata = 32'd64292;
			1245: outdata = 32'd64291;
			1246: outdata = 32'd64290;
			1247: outdata = 32'd64289;
			1248: outdata = 32'd64288;
			1249: outdata = 32'd64287;
			1250: outdata = 32'd64286;
			1251: outdata = 32'd64285;
			1252: outdata = 32'd64284;
			1253: outdata = 32'd64283;
			1254: outdata = 32'd64282;
			1255: outdata = 32'd64281;
			1256: outdata = 32'd64280;
			1257: outdata = 32'd64279;
			1258: outdata = 32'd64278;
			1259: outdata = 32'd64277;
			1260: outdata = 32'd64276;
			1261: outdata = 32'd64275;
			1262: outdata = 32'd64274;
			1263: outdata = 32'd64273;
			1264: outdata = 32'd64272;
			1265: outdata = 32'd64271;
			1266: outdata = 32'd64270;
			1267: outdata = 32'd64269;
			1268: outdata = 32'd64268;
			1269: outdata = 32'd64267;
			1270: outdata = 32'd64266;
			1271: outdata = 32'd64265;
			1272: outdata = 32'd64264;
			1273: outdata = 32'd64263;
			1274: outdata = 32'd64262;
			1275: outdata = 32'd64261;
			1276: outdata = 32'd64260;
			1277: outdata = 32'd64259;
			1278: outdata = 32'd64258;
			1279: outdata = 32'd64257;
			1280: outdata = 32'd64256;
			1281: outdata = 32'd64255;
			1282: outdata = 32'd64254;
			1283: outdata = 32'd64253;
			1284: outdata = 32'd64252;
			1285: outdata = 32'd64251;
			1286: outdata = 32'd64250;
			1287: outdata = 32'd64249;
			1288: outdata = 32'd64248;
			1289: outdata = 32'd64247;
			1290: outdata = 32'd64246;
			1291: outdata = 32'd64245;
			1292: outdata = 32'd64244;
			1293: outdata = 32'd64243;
			1294: outdata = 32'd64242;
			1295: outdata = 32'd64241;
			1296: outdata = 32'd64240;
			1297: outdata = 32'd64239;
			1298: outdata = 32'd64238;
			1299: outdata = 32'd64237;
			1300: outdata = 32'd64236;
			1301: outdata = 32'd64235;
			1302: outdata = 32'd64234;
			1303: outdata = 32'd64233;
			1304: outdata = 32'd64232;
			1305: outdata = 32'd64231;
			1306: outdata = 32'd64230;
			1307: outdata = 32'd64229;
			1308: outdata = 32'd64228;
			1309: outdata = 32'd64227;
			1310: outdata = 32'd64226;
			1311: outdata = 32'd64225;
			1312: outdata = 32'd64224;
			1313: outdata = 32'd64223;
			1314: outdata = 32'd64222;
			1315: outdata = 32'd64221;
			1316: outdata = 32'd64220;
			1317: outdata = 32'd64219;
			1318: outdata = 32'd64218;
			1319: outdata = 32'd64217;
			1320: outdata = 32'd64216;
			1321: outdata = 32'd64215;
			1322: outdata = 32'd64214;
			1323: outdata = 32'd64213;
			1324: outdata = 32'd64212;
			1325: outdata = 32'd64211;
			1326: outdata = 32'd64210;
			1327: outdata = 32'd64209;
			1328: outdata = 32'd64208;
			1329: outdata = 32'd64207;
			1330: outdata = 32'd64206;
			1331: outdata = 32'd64205;
			1332: outdata = 32'd64204;
			1333: outdata = 32'd64203;
			1334: outdata = 32'd64202;
			1335: outdata = 32'd64201;
			1336: outdata = 32'd64200;
			1337: outdata = 32'd64199;
			1338: outdata = 32'd64198;
			1339: outdata = 32'd64197;
			1340: outdata = 32'd64196;
			1341: outdata = 32'd64195;
			1342: outdata = 32'd64194;
			1343: outdata = 32'd64193;
			1344: outdata = 32'd64192;
			1345: outdata = 32'd64191;
			1346: outdata = 32'd64190;
			1347: outdata = 32'd64189;
			1348: outdata = 32'd64188;
			1349: outdata = 32'd64187;
			1350: outdata = 32'd64186;
			1351: outdata = 32'd64185;
			1352: outdata = 32'd64184;
			1353: outdata = 32'd64183;
			1354: outdata = 32'd64182;
			1355: outdata = 32'd64181;
			1356: outdata = 32'd64180;
			1357: outdata = 32'd64179;
			1358: outdata = 32'd64178;
			1359: outdata = 32'd64177;
			1360: outdata = 32'd64176;
			1361: outdata = 32'd64175;
			1362: outdata = 32'd64174;
			1363: outdata = 32'd64173;
			1364: outdata = 32'd64172;
			1365: outdata = 32'd64171;
			1366: outdata = 32'd64170;
			1367: outdata = 32'd64169;
			1368: outdata = 32'd64168;
			1369: outdata = 32'd64167;
			1370: outdata = 32'd64166;
			1371: outdata = 32'd64165;
			1372: outdata = 32'd64164;
			1373: outdata = 32'd64163;
			1374: outdata = 32'd64162;
			1375: outdata = 32'd64161;
			1376: outdata = 32'd64160;
			1377: outdata = 32'd64159;
			1378: outdata = 32'd64158;
			1379: outdata = 32'd64157;
			1380: outdata = 32'd64156;
			1381: outdata = 32'd64155;
			1382: outdata = 32'd64154;
			1383: outdata = 32'd64153;
			1384: outdata = 32'd64152;
			1385: outdata = 32'd64151;
			1386: outdata = 32'd64150;
			1387: outdata = 32'd64149;
			1388: outdata = 32'd64148;
			1389: outdata = 32'd64147;
			1390: outdata = 32'd64146;
			1391: outdata = 32'd64145;
			1392: outdata = 32'd64144;
			1393: outdata = 32'd64143;
			1394: outdata = 32'd64142;
			1395: outdata = 32'd64141;
			1396: outdata = 32'd64140;
			1397: outdata = 32'd64139;
			1398: outdata = 32'd64138;
			1399: outdata = 32'd64137;
			1400: outdata = 32'd64136;
			1401: outdata = 32'd64135;
			1402: outdata = 32'd64134;
			1403: outdata = 32'd64133;
			1404: outdata = 32'd64132;
			1405: outdata = 32'd64131;
			1406: outdata = 32'd64130;
			1407: outdata = 32'd64129;
			1408: outdata = 32'd64128;
			1409: outdata = 32'd64127;
			1410: outdata = 32'd64126;
			1411: outdata = 32'd64125;
			1412: outdata = 32'd64124;
			1413: outdata = 32'd64123;
			1414: outdata = 32'd64122;
			1415: outdata = 32'd64121;
			1416: outdata = 32'd64120;
			1417: outdata = 32'd64119;
			1418: outdata = 32'd64118;
			1419: outdata = 32'd64117;
			1420: outdata = 32'd64116;
			1421: outdata = 32'd64115;
			1422: outdata = 32'd64114;
			1423: outdata = 32'd64113;
			1424: outdata = 32'd64112;
			1425: outdata = 32'd64111;
			1426: outdata = 32'd64110;
			1427: outdata = 32'd64109;
			1428: outdata = 32'd64108;
			1429: outdata = 32'd64107;
			1430: outdata = 32'd64106;
			1431: outdata = 32'd64105;
			1432: outdata = 32'd64104;
			1433: outdata = 32'd64103;
			1434: outdata = 32'd64102;
			1435: outdata = 32'd64101;
			1436: outdata = 32'd64100;
			1437: outdata = 32'd64099;
			1438: outdata = 32'd64098;
			1439: outdata = 32'd64097;
			1440: outdata = 32'd64096;
			1441: outdata = 32'd64095;
			1442: outdata = 32'd64094;
			1443: outdata = 32'd64093;
			1444: outdata = 32'd64092;
			1445: outdata = 32'd64091;
			1446: outdata = 32'd64090;
			1447: outdata = 32'd64089;
			1448: outdata = 32'd64088;
			1449: outdata = 32'd64087;
			1450: outdata = 32'd64086;
			1451: outdata = 32'd64085;
			1452: outdata = 32'd64084;
			1453: outdata = 32'd64083;
			1454: outdata = 32'd64082;
			1455: outdata = 32'd64081;
			1456: outdata = 32'd64080;
			1457: outdata = 32'd64079;
			1458: outdata = 32'd64078;
			1459: outdata = 32'd64077;
			1460: outdata = 32'd64076;
			1461: outdata = 32'd64075;
			1462: outdata = 32'd64074;
			1463: outdata = 32'd64073;
			1464: outdata = 32'd64072;
			1465: outdata = 32'd64071;
			1466: outdata = 32'd64070;
			1467: outdata = 32'd64069;
			1468: outdata = 32'd64068;
			1469: outdata = 32'd64067;
			1470: outdata = 32'd64066;
			1471: outdata = 32'd64065;
			1472: outdata = 32'd64064;
			1473: outdata = 32'd64063;
			1474: outdata = 32'd64062;
			1475: outdata = 32'd64061;
			1476: outdata = 32'd64060;
			1477: outdata = 32'd64059;
			1478: outdata = 32'd64058;
			1479: outdata = 32'd64057;
			1480: outdata = 32'd64056;
			1481: outdata = 32'd64055;
			1482: outdata = 32'd64054;
			1483: outdata = 32'd64053;
			1484: outdata = 32'd64052;
			1485: outdata = 32'd64051;
			1486: outdata = 32'd64050;
			1487: outdata = 32'd64049;
			1488: outdata = 32'd64048;
			1489: outdata = 32'd64047;
			1490: outdata = 32'd64046;
			1491: outdata = 32'd64045;
			1492: outdata = 32'd64044;
			1493: outdata = 32'd64043;
			1494: outdata = 32'd64042;
			1495: outdata = 32'd64041;
			1496: outdata = 32'd64040;
			1497: outdata = 32'd64039;
			1498: outdata = 32'd64038;
			1499: outdata = 32'd64037;
			1500: outdata = 32'd64036;
			1501: outdata = 32'd64035;
			1502: outdata = 32'd64034;
			1503: outdata = 32'd64033;
			1504: outdata = 32'd64032;
			1505: outdata = 32'd64031;
			1506: outdata = 32'd64030;
			1507: outdata = 32'd64029;
			1508: outdata = 32'd64028;
			1509: outdata = 32'd64027;
			1510: outdata = 32'd64026;
			1511: outdata = 32'd64025;
			1512: outdata = 32'd64024;
			1513: outdata = 32'd64023;
			1514: outdata = 32'd64022;
			1515: outdata = 32'd64021;
			1516: outdata = 32'd64020;
			1517: outdata = 32'd64019;
			1518: outdata = 32'd64018;
			1519: outdata = 32'd64017;
			1520: outdata = 32'd64016;
			1521: outdata = 32'd64015;
			1522: outdata = 32'd64014;
			1523: outdata = 32'd64013;
			1524: outdata = 32'd64012;
			1525: outdata = 32'd64011;
			1526: outdata = 32'd64010;
			1527: outdata = 32'd64009;
			1528: outdata = 32'd64008;
			1529: outdata = 32'd64007;
			1530: outdata = 32'd64006;
			1531: outdata = 32'd64005;
			1532: outdata = 32'd64004;
			1533: outdata = 32'd64003;
			1534: outdata = 32'd64002;
			1535: outdata = 32'd64001;
			1536: outdata = 32'd64000;
			1537: outdata = 32'd63999;
			1538: outdata = 32'd63998;
			1539: outdata = 32'd63997;
			1540: outdata = 32'd63996;
			1541: outdata = 32'd63995;
			1542: outdata = 32'd63994;
			1543: outdata = 32'd63993;
			1544: outdata = 32'd63992;
			1545: outdata = 32'd63991;
			1546: outdata = 32'd63990;
			1547: outdata = 32'd63989;
			1548: outdata = 32'd63988;
			1549: outdata = 32'd63987;
			1550: outdata = 32'd63986;
			1551: outdata = 32'd63985;
			1552: outdata = 32'd63984;
			1553: outdata = 32'd63983;
			1554: outdata = 32'd63982;
			1555: outdata = 32'd63981;
			1556: outdata = 32'd63980;
			1557: outdata = 32'd63979;
			1558: outdata = 32'd63978;
			1559: outdata = 32'd63977;
			1560: outdata = 32'd63976;
			1561: outdata = 32'd63975;
			1562: outdata = 32'd63974;
			1563: outdata = 32'd63973;
			1564: outdata = 32'd63972;
			1565: outdata = 32'd63971;
			1566: outdata = 32'd63970;
			1567: outdata = 32'd63969;
			1568: outdata = 32'd63968;
			1569: outdata = 32'd63967;
			1570: outdata = 32'd63966;
			1571: outdata = 32'd63965;
			1572: outdata = 32'd63964;
			1573: outdata = 32'd63963;
			1574: outdata = 32'd63962;
			1575: outdata = 32'd63961;
			1576: outdata = 32'd63960;
			1577: outdata = 32'd63959;
			1578: outdata = 32'd63958;
			1579: outdata = 32'd63957;
			1580: outdata = 32'd63956;
			1581: outdata = 32'd63955;
			1582: outdata = 32'd63954;
			1583: outdata = 32'd63953;
			1584: outdata = 32'd63952;
			1585: outdata = 32'd63951;
			1586: outdata = 32'd63950;
			1587: outdata = 32'd63949;
			1588: outdata = 32'd63948;
			1589: outdata = 32'd63947;
			1590: outdata = 32'd63946;
			1591: outdata = 32'd63945;
			1592: outdata = 32'd63944;
			1593: outdata = 32'd63943;
			1594: outdata = 32'd63942;
			1595: outdata = 32'd63941;
			1596: outdata = 32'd63940;
			1597: outdata = 32'd63939;
			1598: outdata = 32'd63938;
			1599: outdata = 32'd63937;
			1600: outdata = 32'd63936;
			1601: outdata = 32'd63935;
			1602: outdata = 32'd63934;
			1603: outdata = 32'd63933;
			1604: outdata = 32'd63932;
			1605: outdata = 32'd63931;
			1606: outdata = 32'd63930;
			1607: outdata = 32'd63929;
			1608: outdata = 32'd63928;
			1609: outdata = 32'd63927;
			1610: outdata = 32'd63926;
			1611: outdata = 32'd63925;
			1612: outdata = 32'd63924;
			1613: outdata = 32'd63923;
			1614: outdata = 32'd63922;
			1615: outdata = 32'd63921;
			1616: outdata = 32'd63920;
			1617: outdata = 32'd63919;
			1618: outdata = 32'd63918;
			1619: outdata = 32'd63917;
			1620: outdata = 32'd63916;
			1621: outdata = 32'd63915;
			1622: outdata = 32'd63914;
			1623: outdata = 32'd63913;
			1624: outdata = 32'd63912;
			1625: outdata = 32'd63911;
			1626: outdata = 32'd63910;
			1627: outdata = 32'd63909;
			1628: outdata = 32'd63908;
			1629: outdata = 32'd63907;
			1630: outdata = 32'd63906;
			1631: outdata = 32'd63905;
			1632: outdata = 32'd63904;
			1633: outdata = 32'd63903;
			1634: outdata = 32'd63902;
			1635: outdata = 32'd63901;
			1636: outdata = 32'd63900;
			1637: outdata = 32'd63899;
			1638: outdata = 32'd63898;
			1639: outdata = 32'd63897;
			1640: outdata = 32'd63896;
			1641: outdata = 32'd63895;
			1642: outdata = 32'd63894;
			1643: outdata = 32'd63893;
			1644: outdata = 32'd63892;
			1645: outdata = 32'd63891;
			1646: outdata = 32'd63890;
			1647: outdata = 32'd63889;
			1648: outdata = 32'd63888;
			1649: outdata = 32'd63887;
			1650: outdata = 32'd63886;
			1651: outdata = 32'd63885;
			1652: outdata = 32'd63884;
			1653: outdata = 32'd63883;
			1654: outdata = 32'd63882;
			1655: outdata = 32'd63881;
			1656: outdata = 32'd63880;
			1657: outdata = 32'd63879;
			1658: outdata = 32'd63878;
			1659: outdata = 32'd63877;
			1660: outdata = 32'd63876;
			1661: outdata = 32'd63875;
			1662: outdata = 32'd63874;
			1663: outdata = 32'd63873;
			1664: outdata = 32'd63872;
			1665: outdata = 32'd63871;
			1666: outdata = 32'd63870;
			1667: outdata = 32'd63869;
			1668: outdata = 32'd63868;
			1669: outdata = 32'd63867;
			1670: outdata = 32'd63866;
			1671: outdata = 32'd63865;
			1672: outdata = 32'd63864;
			1673: outdata = 32'd63863;
			1674: outdata = 32'd63862;
			1675: outdata = 32'd63861;
			1676: outdata = 32'd63860;
			1677: outdata = 32'd63859;
			1678: outdata = 32'd63858;
			1679: outdata = 32'd63857;
			1680: outdata = 32'd63856;
			1681: outdata = 32'd63855;
			1682: outdata = 32'd63854;
			1683: outdata = 32'd63853;
			1684: outdata = 32'd63852;
			1685: outdata = 32'd63851;
			1686: outdata = 32'd63850;
			1687: outdata = 32'd63849;
			1688: outdata = 32'd63848;
			1689: outdata = 32'd63847;
			1690: outdata = 32'd63846;
			1691: outdata = 32'd63845;
			1692: outdata = 32'd63844;
			1693: outdata = 32'd63843;
			1694: outdata = 32'd63842;
			1695: outdata = 32'd63841;
			1696: outdata = 32'd63840;
			1697: outdata = 32'd63839;
			1698: outdata = 32'd63838;
			1699: outdata = 32'd63837;
			1700: outdata = 32'd63836;
			1701: outdata = 32'd63835;
			1702: outdata = 32'd63834;
			1703: outdata = 32'd63833;
			1704: outdata = 32'd63832;
			1705: outdata = 32'd63831;
			1706: outdata = 32'd63830;
			1707: outdata = 32'd63829;
			1708: outdata = 32'd63828;
			1709: outdata = 32'd63827;
			1710: outdata = 32'd63826;
			1711: outdata = 32'd63825;
			1712: outdata = 32'd63824;
			1713: outdata = 32'd63823;
			1714: outdata = 32'd63822;
			1715: outdata = 32'd63821;
			1716: outdata = 32'd63820;
			1717: outdata = 32'd63819;
			1718: outdata = 32'd63818;
			1719: outdata = 32'd63817;
			1720: outdata = 32'd63816;
			1721: outdata = 32'd63815;
			1722: outdata = 32'd63814;
			1723: outdata = 32'd63813;
			1724: outdata = 32'd63812;
			1725: outdata = 32'd63811;
			1726: outdata = 32'd63810;
			1727: outdata = 32'd63809;
			1728: outdata = 32'd63808;
			1729: outdata = 32'd63807;
			1730: outdata = 32'd63806;
			1731: outdata = 32'd63805;
			1732: outdata = 32'd63804;
			1733: outdata = 32'd63803;
			1734: outdata = 32'd63802;
			1735: outdata = 32'd63801;
			1736: outdata = 32'd63800;
			1737: outdata = 32'd63799;
			1738: outdata = 32'd63798;
			1739: outdata = 32'd63797;
			1740: outdata = 32'd63796;
			1741: outdata = 32'd63795;
			1742: outdata = 32'd63794;
			1743: outdata = 32'd63793;
			1744: outdata = 32'd63792;
			1745: outdata = 32'd63791;
			1746: outdata = 32'd63790;
			1747: outdata = 32'd63789;
			1748: outdata = 32'd63788;
			1749: outdata = 32'd63787;
			1750: outdata = 32'd63786;
			1751: outdata = 32'd63785;
			1752: outdata = 32'd63784;
			1753: outdata = 32'd63783;
			1754: outdata = 32'd63782;
			1755: outdata = 32'd63781;
			1756: outdata = 32'd63780;
			1757: outdata = 32'd63779;
			1758: outdata = 32'd63778;
			1759: outdata = 32'd63777;
			1760: outdata = 32'd63776;
			1761: outdata = 32'd63775;
			1762: outdata = 32'd63774;
			1763: outdata = 32'd63773;
			1764: outdata = 32'd63772;
			1765: outdata = 32'd63771;
			1766: outdata = 32'd63770;
			1767: outdata = 32'd63769;
			1768: outdata = 32'd63768;
			1769: outdata = 32'd63767;
			1770: outdata = 32'd63766;
			1771: outdata = 32'd63765;
			1772: outdata = 32'd63764;
			1773: outdata = 32'd63763;
			1774: outdata = 32'd63762;
			1775: outdata = 32'd63761;
			1776: outdata = 32'd63760;
			1777: outdata = 32'd63759;
			1778: outdata = 32'd63758;
			1779: outdata = 32'd63757;
			1780: outdata = 32'd63756;
			1781: outdata = 32'd63755;
			1782: outdata = 32'd63754;
			1783: outdata = 32'd63753;
			1784: outdata = 32'd63752;
			1785: outdata = 32'd63751;
			1786: outdata = 32'd63750;
			1787: outdata = 32'd63749;
			1788: outdata = 32'd63748;
			1789: outdata = 32'd63747;
			1790: outdata = 32'd63746;
			1791: outdata = 32'd63745;
			1792: outdata = 32'd63744;
			1793: outdata = 32'd63743;
			1794: outdata = 32'd63742;
			1795: outdata = 32'd63741;
			1796: outdata = 32'd63740;
			1797: outdata = 32'd63739;
			1798: outdata = 32'd63738;
			1799: outdata = 32'd63737;
			1800: outdata = 32'd63736;
			1801: outdata = 32'd63735;
			1802: outdata = 32'd63734;
			1803: outdata = 32'd63733;
			1804: outdata = 32'd63732;
			1805: outdata = 32'd63731;
			1806: outdata = 32'd63730;
			1807: outdata = 32'd63729;
			1808: outdata = 32'd63728;
			1809: outdata = 32'd63727;
			1810: outdata = 32'd63726;
			1811: outdata = 32'd63725;
			1812: outdata = 32'd63724;
			1813: outdata = 32'd63723;
			1814: outdata = 32'd63722;
			1815: outdata = 32'd63721;
			1816: outdata = 32'd63720;
			1817: outdata = 32'd63719;
			1818: outdata = 32'd63718;
			1819: outdata = 32'd63717;
			1820: outdata = 32'd63716;
			1821: outdata = 32'd63715;
			1822: outdata = 32'd63714;
			1823: outdata = 32'd63713;
			1824: outdata = 32'd63712;
			1825: outdata = 32'd63711;
			1826: outdata = 32'd63710;
			1827: outdata = 32'd63709;
			1828: outdata = 32'd63708;
			1829: outdata = 32'd63707;
			1830: outdata = 32'd63706;
			1831: outdata = 32'd63705;
			1832: outdata = 32'd63704;
			1833: outdata = 32'd63703;
			1834: outdata = 32'd63702;
			1835: outdata = 32'd63701;
			1836: outdata = 32'd63700;
			1837: outdata = 32'd63699;
			1838: outdata = 32'd63698;
			1839: outdata = 32'd63697;
			1840: outdata = 32'd63696;
			1841: outdata = 32'd63695;
			1842: outdata = 32'd63694;
			1843: outdata = 32'd63693;
			1844: outdata = 32'd63692;
			1845: outdata = 32'd63691;
			1846: outdata = 32'd63690;
			1847: outdata = 32'd63689;
			1848: outdata = 32'd63688;
			1849: outdata = 32'd63687;
			1850: outdata = 32'd63686;
			1851: outdata = 32'd63685;
			1852: outdata = 32'd63684;
			1853: outdata = 32'd63683;
			1854: outdata = 32'd63682;
			1855: outdata = 32'd63681;
			1856: outdata = 32'd63680;
			1857: outdata = 32'd63679;
			1858: outdata = 32'd63678;
			1859: outdata = 32'd63677;
			1860: outdata = 32'd63676;
			1861: outdata = 32'd63675;
			1862: outdata = 32'd63674;
			1863: outdata = 32'd63673;
			1864: outdata = 32'd63672;
			1865: outdata = 32'd63671;
			1866: outdata = 32'd63670;
			1867: outdata = 32'd63669;
			1868: outdata = 32'd63668;
			1869: outdata = 32'd63667;
			1870: outdata = 32'd63666;
			1871: outdata = 32'd63665;
			1872: outdata = 32'd63664;
			1873: outdata = 32'd63663;
			1874: outdata = 32'd63662;
			1875: outdata = 32'd63661;
			1876: outdata = 32'd63660;
			1877: outdata = 32'd63659;
			1878: outdata = 32'd63658;
			1879: outdata = 32'd63657;
			1880: outdata = 32'd63656;
			1881: outdata = 32'd63655;
			1882: outdata = 32'd63654;
			1883: outdata = 32'd63653;
			1884: outdata = 32'd63652;
			1885: outdata = 32'd63651;
			1886: outdata = 32'd63650;
			1887: outdata = 32'd63649;
			1888: outdata = 32'd63648;
			1889: outdata = 32'd63647;
			1890: outdata = 32'd63646;
			1891: outdata = 32'd63645;
			1892: outdata = 32'd63644;
			1893: outdata = 32'd63643;
			1894: outdata = 32'd63642;
			1895: outdata = 32'd63641;
			1896: outdata = 32'd63640;
			1897: outdata = 32'd63639;
			1898: outdata = 32'd63638;
			1899: outdata = 32'd63637;
			1900: outdata = 32'd63636;
			1901: outdata = 32'd63635;
			1902: outdata = 32'd63634;
			1903: outdata = 32'd63633;
			1904: outdata = 32'd63632;
			1905: outdata = 32'd63631;
			1906: outdata = 32'd63630;
			1907: outdata = 32'd63629;
			1908: outdata = 32'd63628;
			1909: outdata = 32'd63627;
			1910: outdata = 32'd63626;
			1911: outdata = 32'd63625;
			1912: outdata = 32'd63624;
			1913: outdata = 32'd63623;
			1914: outdata = 32'd63622;
			1915: outdata = 32'd63621;
			1916: outdata = 32'd63620;
			1917: outdata = 32'd63619;
			1918: outdata = 32'd63618;
			1919: outdata = 32'd63617;
			1920: outdata = 32'd63616;
			1921: outdata = 32'd63615;
			1922: outdata = 32'd63614;
			1923: outdata = 32'd63613;
			1924: outdata = 32'd63612;
			1925: outdata = 32'd63611;
			1926: outdata = 32'd63610;
			1927: outdata = 32'd63609;
			1928: outdata = 32'd63608;
			1929: outdata = 32'd63607;
			1930: outdata = 32'd63606;
			1931: outdata = 32'd63605;
			1932: outdata = 32'd63604;
			1933: outdata = 32'd63603;
			1934: outdata = 32'd63602;
			1935: outdata = 32'd63601;
			1936: outdata = 32'd63600;
			1937: outdata = 32'd63599;
			1938: outdata = 32'd63598;
			1939: outdata = 32'd63597;
			1940: outdata = 32'd63596;
			1941: outdata = 32'd63595;
			1942: outdata = 32'd63594;
			1943: outdata = 32'd63593;
			1944: outdata = 32'd63592;
			1945: outdata = 32'd63591;
			1946: outdata = 32'd63590;
			1947: outdata = 32'd63589;
			1948: outdata = 32'd63588;
			1949: outdata = 32'd63587;
			1950: outdata = 32'd63586;
			1951: outdata = 32'd63585;
			1952: outdata = 32'd63584;
			1953: outdata = 32'd63583;
			1954: outdata = 32'd63582;
			1955: outdata = 32'd63581;
			1956: outdata = 32'd63580;
			1957: outdata = 32'd63579;
			1958: outdata = 32'd63578;
			1959: outdata = 32'd63577;
			1960: outdata = 32'd63576;
			1961: outdata = 32'd63575;
			1962: outdata = 32'd63574;
			1963: outdata = 32'd63573;
			1964: outdata = 32'd63572;
			1965: outdata = 32'd63571;
			1966: outdata = 32'd63570;
			1967: outdata = 32'd63569;
			1968: outdata = 32'd63568;
			1969: outdata = 32'd63567;
			1970: outdata = 32'd63566;
			1971: outdata = 32'd63565;
			1972: outdata = 32'd63564;
			1973: outdata = 32'd63563;
			1974: outdata = 32'd63562;
			1975: outdata = 32'd63561;
			1976: outdata = 32'd63560;
			1977: outdata = 32'd63559;
			1978: outdata = 32'd63558;
			1979: outdata = 32'd63557;
			1980: outdata = 32'd63556;
			1981: outdata = 32'd63555;
			1982: outdata = 32'd63554;
			1983: outdata = 32'd63553;
			1984: outdata = 32'd63552;
			1985: outdata = 32'd63551;
			1986: outdata = 32'd63550;
			1987: outdata = 32'd63549;
			1988: outdata = 32'd63548;
			1989: outdata = 32'd63547;
			1990: outdata = 32'd63546;
			1991: outdata = 32'd63545;
			1992: outdata = 32'd63544;
			1993: outdata = 32'd63543;
			1994: outdata = 32'd63542;
			1995: outdata = 32'd63541;
			1996: outdata = 32'd63540;
			1997: outdata = 32'd63539;
			1998: outdata = 32'd63538;
			1999: outdata = 32'd63537;
			2000: outdata = 32'd63536;
			2001: outdata = 32'd63535;
			2002: outdata = 32'd63534;
			2003: outdata = 32'd63533;
			2004: outdata = 32'd63532;
			2005: outdata = 32'd63531;
			2006: outdata = 32'd63530;
			2007: outdata = 32'd63529;
			2008: outdata = 32'd63528;
			2009: outdata = 32'd63527;
			2010: outdata = 32'd63526;
			2011: outdata = 32'd63525;
			2012: outdata = 32'd63524;
			2013: outdata = 32'd63523;
			2014: outdata = 32'd63522;
			2015: outdata = 32'd63521;
			2016: outdata = 32'd63520;
			2017: outdata = 32'd63519;
			2018: outdata = 32'd63518;
			2019: outdata = 32'd63517;
			2020: outdata = 32'd63516;
			2021: outdata = 32'd63515;
			2022: outdata = 32'd63514;
			2023: outdata = 32'd63513;
			2024: outdata = 32'd63512;
			2025: outdata = 32'd63511;
			2026: outdata = 32'd63510;
			2027: outdata = 32'd63509;
			2028: outdata = 32'd63508;
			2029: outdata = 32'd63507;
			2030: outdata = 32'd63506;
			2031: outdata = 32'd63505;
			2032: outdata = 32'd63504;
			2033: outdata = 32'd63503;
			2034: outdata = 32'd63502;
			2035: outdata = 32'd63501;
			2036: outdata = 32'd63500;
			2037: outdata = 32'd63499;
			2038: outdata = 32'd63498;
			2039: outdata = 32'd63497;
			2040: outdata = 32'd63496;
			2041: outdata = 32'd63495;
			2042: outdata = 32'd63494;
			2043: outdata = 32'd63493;
			2044: outdata = 32'd63492;
			2045: outdata = 32'd63491;
			2046: outdata = 32'd63490;
			2047: outdata = 32'd63489;
			2048: outdata = 32'd63488;
			2049: outdata = 32'd63487;
			2050: outdata = 32'd63486;
			2051: outdata = 32'd63485;
			2052: outdata = 32'd63484;
			2053: outdata = 32'd63483;
			2054: outdata = 32'd63482;
			2055: outdata = 32'd63481;
			2056: outdata = 32'd63480;
			2057: outdata = 32'd63479;
			2058: outdata = 32'd63478;
			2059: outdata = 32'd63477;
			2060: outdata = 32'd63476;
			2061: outdata = 32'd63475;
			2062: outdata = 32'd63474;
			2063: outdata = 32'd63473;
			2064: outdata = 32'd63472;
			2065: outdata = 32'd63471;
			2066: outdata = 32'd63470;
			2067: outdata = 32'd63469;
			2068: outdata = 32'd63468;
			2069: outdata = 32'd63467;
			2070: outdata = 32'd63466;
			2071: outdata = 32'd63465;
			2072: outdata = 32'd63464;
			2073: outdata = 32'd63463;
			2074: outdata = 32'd63462;
			2075: outdata = 32'd63461;
			2076: outdata = 32'd63460;
			2077: outdata = 32'd63459;
			2078: outdata = 32'd63458;
			2079: outdata = 32'd63457;
			2080: outdata = 32'd63456;
			2081: outdata = 32'd63455;
			2082: outdata = 32'd63454;
			2083: outdata = 32'd63453;
			2084: outdata = 32'd63452;
			2085: outdata = 32'd63451;
			2086: outdata = 32'd63450;
			2087: outdata = 32'd63449;
			2088: outdata = 32'd63448;
			2089: outdata = 32'd63447;
			2090: outdata = 32'd63446;
			2091: outdata = 32'd63445;
			2092: outdata = 32'd63444;
			2093: outdata = 32'd63443;
			2094: outdata = 32'd63442;
			2095: outdata = 32'd63441;
			2096: outdata = 32'd63440;
			2097: outdata = 32'd63439;
			2098: outdata = 32'd63438;
			2099: outdata = 32'd63437;
			2100: outdata = 32'd63436;
			2101: outdata = 32'd63435;
			2102: outdata = 32'd63434;
			2103: outdata = 32'd63433;
			2104: outdata = 32'd63432;
			2105: outdata = 32'd63431;
			2106: outdata = 32'd63430;
			2107: outdata = 32'd63429;
			2108: outdata = 32'd63428;
			2109: outdata = 32'd63427;
			2110: outdata = 32'd63426;
			2111: outdata = 32'd63425;
			2112: outdata = 32'd63424;
			2113: outdata = 32'd63423;
			2114: outdata = 32'd63422;
			2115: outdata = 32'd63421;
			2116: outdata = 32'd63420;
			2117: outdata = 32'd63419;
			2118: outdata = 32'd63418;
			2119: outdata = 32'd63417;
			2120: outdata = 32'd63416;
			2121: outdata = 32'd63415;
			2122: outdata = 32'd63414;
			2123: outdata = 32'd63413;
			2124: outdata = 32'd63412;
			2125: outdata = 32'd63411;
			2126: outdata = 32'd63410;
			2127: outdata = 32'd63409;
			2128: outdata = 32'd63408;
			2129: outdata = 32'd63407;
			2130: outdata = 32'd63406;
			2131: outdata = 32'd63405;
			2132: outdata = 32'd63404;
			2133: outdata = 32'd63403;
			2134: outdata = 32'd63402;
			2135: outdata = 32'd63401;
			2136: outdata = 32'd63400;
			2137: outdata = 32'd63399;
			2138: outdata = 32'd63398;
			2139: outdata = 32'd63397;
			2140: outdata = 32'd63396;
			2141: outdata = 32'd63395;
			2142: outdata = 32'd63394;
			2143: outdata = 32'd63393;
			2144: outdata = 32'd63392;
			2145: outdata = 32'd63391;
			2146: outdata = 32'd63390;
			2147: outdata = 32'd63389;
			2148: outdata = 32'd63388;
			2149: outdata = 32'd63387;
			2150: outdata = 32'd63386;
			2151: outdata = 32'd63385;
			2152: outdata = 32'd63384;
			2153: outdata = 32'd63383;
			2154: outdata = 32'd63382;
			2155: outdata = 32'd63381;
			2156: outdata = 32'd63380;
			2157: outdata = 32'd63379;
			2158: outdata = 32'd63378;
			2159: outdata = 32'd63377;
			2160: outdata = 32'd63376;
			2161: outdata = 32'd63375;
			2162: outdata = 32'd63374;
			2163: outdata = 32'd63373;
			2164: outdata = 32'd63372;
			2165: outdata = 32'd63371;
			2166: outdata = 32'd63370;
			2167: outdata = 32'd63369;
			2168: outdata = 32'd63368;
			2169: outdata = 32'd63367;
			2170: outdata = 32'd63366;
			2171: outdata = 32'd63365;
			2172: outdata = 32'd63364;
			2173: outdata = 32'd63363;
			2174: outdata = 32'd63362;
			2175: outdata = 32'd63361;
			2176: outdata = 32'd63360;
			2177: outdata = 32'd63359;
			2178: outdata = 32'd63358;
			2179: outdata = 32'd63357;
			2180: outdata = 32'd63356;
			2181: outdata = 32'd63355;
			2182: outdata = 32'd63354;
			2183: outdata = 32'd63353;
			2184: outdata = 32'd63352;
			2185: outdata = 32'd63351;
			2186: outdata = 32'd63350;
			2187: outdata = 32'd63349;
			2188: outdata = 32'd63348;
			2189: outdata = 32'd63347;
			2190: outdata = 32'd63346;
			2191: outdata = 32'd63345;
			2192: outdata = 32'd63344;
			2193: outdata = 32'd63343;
			2194: outdata = 32'd63342;
			2195: outdata = 32'd63341;
			2196: outdata = 32'd63340;
			2197: outdata = 32'd63339;
			2198: outdata = 32'd63338;
			2199: outdata = 32'd63337;
			2200: outdata = 32'd63336;
			2201: outdata = 32'd63335;
			2202: outdata = 32'd63334;
			2203: outdata = 32'd63333;
			2204: outdata = 32'd63332;
			2205: outdata = 32'd63331;
			2206: outdata = 32'd63330;
			2207: outdata = 32'd63329;
			2208: outdata = 32'd63328;
			2209: outdata = 32'd63327;
			2210: outdata = 32'd63326;
			2211: outdata = 32'd63325;
			2212: outdata = 32'd63324;
			2213: outdata = 32'd63323;
			2214: outdata = 32'd63322;
			2215: outdata = 32'd63321;
			2216: outdata = 32'd63320;
			2217: outdata = 32'd63319;
			2218: outdata = 32'd63318;
			2219: outdata = 32'd63317;
			2220: outdata = 32'd63316;
			2221: outdata = 32'd63315;
			2222: outdata = 32'd63314;
			2223: outdata = 32'd63313;
			2224: outdata = 32'd63312;
			2225: outdata = 32'd63311;
			2226: outdata = 32'd63310;
			2227: outdata = 32'd63309;
			2228: outdata = 32'd63308;
			2229: outdata = 32'd63307;
			2230: outdata = 32'd63306;
			2231: outdata = 32'd63305;
			2232: outdata = 32'd63304;
			2233: outdata = 32'd63303;
			2234: outdata = 32'd63302;
			2235: outdata = 32'd63301;
			2236: outdata = 32'd63300;
			2237: outdata = 32'd63299;
			2238: outdata = 32'd63298;
			2239: outdata = 32'd63297;
			2240: outdata = 32'd63296;
			2241: outdata = 32'd63295;
			2242: outdata = 32'd63294;
			2243: outdata = 32'd63293;
			2244: outdata = 32'd63292;
			2245: outdata = 32'd63291;
			2246: outdata = 32'd63290;
			2247: outdata = 32'd63289;
			2248: outdata = 32'd63288;
			2249: outdata = 32'd63287;
			2250: outdata = 32'd63286;
			2251: outdata = 32'd63285;
			2252: outdata = 32'd63284;
			2253: outdata = 32'd63283;
			2254: outdata = 32'd63282;
			2255: outdata = 32'd63281;
			2256: outdata = 32'd63280;
			2257: outdata = 32'd63279;
			2258: outdata = 32'd63278;
			2259: outdata = 32'd63277;
			2260: outdata = 32'd63276;
			2261: outdata = 32'd63275;
			2262: outdata = 32'd63274;
			2263: outdata = 32'd63273;
			2264: outdata = 32'd63272;
			2265: outdata = 32'd63271;
			2266: outdata = 32'd63270;
			2267: outdata = 32'd63269;
			2268: outdata = 32'd63268;
			2269: outdata = 32'd63267;
			2270: outdata = 32'd63266;
			2271: outdata = 32'd63265;
			2272: outdata = 32'd63264;
			2273: outdata = 32'd63263;
			2274: outdata = 32'd63262;
			2275: outdata = 32'd63261;
			2276: outdata = 32'd63260;
			2277: outdata = 32'd63259;
			2278: outdata = 32'd63258;
			2279: outdata = 32'd63257;
			2280: outdata = 32'd63256;
			2281: outdata = 32'd63255;
			2282: outdata = 32'd63254;
			2283: outdata = 32'd63253;
			2284: outdata = 32'd63252;
			2285: outdata = 32'd63251;
			2286: outdata = 32'd63250;
			2287: outdata = 32'd63249;
			2288: outdata = 32'd63248;
			2289: outdata = 32'd63247;
			2290: outdata = 32'd63246;
			2291: outdata = 32'd63245;
			2292: outdata = 32'd63244;
			2293: outdata = 32'd63243;
			2294: outdata = 32'd63242;
			2295: outdata = 32'd63241;
			2296: outdata = 32'd63240;
			2297: outdata = 32'd63239;
			2298: outdata = 32'd63238;
			2299: outdata = 32'd63237;
			2300: outdata = 32'd63236;
			2301: outdata = 32'd63235;
			2302: outdata = 32'd63234;
			2303: outdata = 32'd63233;
			2304: outdata = 32'd63232;
			2305: outdata = 32'd63231;
			2306: outdata = 32'd63230;
			2307: outdata = 32'd63229;
			2308: outdata = 32'd63228;
			2309: outdata = 32'd63227;
			2310: outdata = 32'd63226;
			2311: outdata = 32'd63225;
			2312: outdata = 32'd63224;
			2313: outdata = 32'd63223;
			2314: outdata = 32'd63222;
			2315: outdata = 32'd63221;
			2316: outdata = 32'd63220;
			2317: outdata = 32'd63219;
			2318: outdata = 32'd63218;
			2319: outdata = 32'd63217;
			2320: outdata = 32'd63216;
			2321: outdata = 32'd63215;
			2322: outdata = 32'd63214;
			2323: outdata = 32'd63213;
			2324: outdata = 32'd63212;
			2325: outdata = 32'd63211;
			2326: outdata = 32'd63210;
			2327: outdata = 32'd63209;
			2328: outdata = 32'd63208;
			2329: outdata = 32'd63207;
			2330: outdata = 32'd63206;
			2331: outdata = 32'd63205;
			2332: outdata = 32'd63204;
			2333: outdata = 32'd63203;
			2334: outdata = 32'd63202;
			2335: outdata = 32'd63201;
			2336: outdata = 32'd63200;
			2337: outdata = 32'd63199;
			2338: outdata = 32'd63198;
			2339: outdata = 32'd63197;
			2340: outdata = 32'd63196;
			2341: outdata = 32'd63195;
			2342: outdata = 32'd63194;
			2343: outdata = 32'd63193;
			2344: outdata = 32'd63192;
			2345: outdata = 32'd63191;
			2346: outdata = 32'd63190;
			2347: outdata = 32'd63189;
			2348: outdata = 32'd63188;
			2349: outdata = 32'd63187;
			2350: outdata = 32'd63186;
			2351: outdata = 32'd63185;
			2352: outdata = 32'd63184;
			2353: outdata = 32'd63183;
			2354: outdata = 32'd63182;
			2355: outdata = 32'd63181;
			2356: outdata = 32'd63180;
			2357: outdata = 32'd63179;
			2358: outdata = 32'd63178;
			2359: outdata = 32'd63177;
			2360: outdata = 32'd63176;
			2361: outdata = 32'd63175;
			2362: outdata = 32'd63174;
			2363: outdata = 32'd63173;
			2364: outdata = 32'd63172;
			2365: outdata = 32'd63171;
			2366: outdata = 32'd63170;
			2367: outdata = 32'd63169;
			2368: outdata = 32'd63168;
			2369: outdata = 32'd63167;
			2370: outdata = 32'd63166;
			2371: outdata = 32'd63165;
			2372: outdata = 32'd63164;
			2373: outdata = 32'd63163;
			2374: outdata = 32'd63162;
			2375: outdata = 32'd63161;
			2376: outdata = 32'd63160;
			2377: outdata = 32'd63159;
			2378: outdata = 32'd63158;
			2379: outdata = 32'd63157;
			2380: outdata = 32'd63156;
			2381: outdata = 32'd63155;
			2382: outdata = 32'd63154;
			2383: outdata = 32'd63153;
			2384: outdata = 32'd63152;
			2385: outdata = 32'd63151;
			2386: outdata = 32'd63150;
			2387: outdata = 32'd63149;
			2388: outdata = 32'd63148;
			2389: outdata = 32'd63147;
			2390: outdata = 32'd63146;
			2391: outdata = 32'd63145;
			2392: outdata = 32'd63144;
			2393: outdata = 32'd63143;
			2394: outdata = 32'd63142;
			2395: outdata = 32'd63141;
			2396: outdata = 32'd63140;
			2397: outdata = 32'd63139;
			2398: outdata = 32'd63138;
			2399: outdata = 32'd63137;
			2400: outdata = 32'd63136;
			2401: outdata = 32'd63135;
			2402: outdata = 32'd63134;
			2403: outdata = 32'd63133;
			2404: outdata = 32'd63132;
			2405: outdata = 32'd63131;
			2406: outdata = 32'd63130;
			2407: outdata = 32'd63129;
			2408: outdata = 32'd63128;
			2409: outdata = 32'd63127;
			2410: outdata = 32'd63126;
			2411: outdata = 32'd63125;
			2412: outdata = 32'd63124;
			2413: outdata = 32'd63123;
			2414: outdata = 32'd63122;
			2415: outdata = 32'd63121;
			2416: outdata = 32'd63120;
			2417: outdata = 32'd63119;
			2418: outdata = 32'd63118;
			2419: outdata = 32'd63117;
			2420: outdata = 32'd63116;
			2421: outdata = 32'd63115;
			2422: outdata = 32'd63114;
			2423: outdata = 32'd63113;
			2424: outdata = 32'd63112;
			2425: outdata = 32'd63111;
			2426: outdata = 32'd63110;
			2427: outdata = 32'd63109;
			2428: outdata = 32'd63108;
			2429: outdata = 32'd63107;
			2430: outdata = 32'd63106;
			2431: outdata = 32'd63105;
			2432: outdata = 32'd63104;
			2433: outdata = 32'd63103;
			2434: outdata = 32'd63102;
			2435: outdata = 32'd63101;
			2436: outdata = 32'd63100;
			2437: outdata = 32'd63099;
			2438: outdata = 32'd63098;
			2439: outdata = 32'd63097;
			2440: outdata = 32'd63096;
			2441: outdata = 32'd63095;
			2442: outdata = 32'd63094;
			2443: outdata = 32'd63093;
			2444: outdata = 32'd63092;
			2445: outdata = 32'd63091;
			2446: outdata = 32'd63090;
			2447: outdata = 32'd63089;
			2448: outdata = 32'd63088;
			2449: outdata = 32'd63087;
			2450: outdata = 32'd63086;
			2451: outdata = 32'd63085;
			2452: outdata = 32'd63084;
			2453: outdata = 32'd63083;
			2454: outdata = 32'd63082;
			2455: outdata = 32'd63081;
			2456: outdata = 32'd63080;
			2457: outdata = 32'd63079;
			2458: outdata = 32'd63078;
			2459: outdata = 32'd63077;
			2460: outdata = 32'd63076;
			2461: outdata = 32'd63075;
			2462: outdata = 32'd63074;
			2463: outdata = 32'd63073;
			2464: outdata = 32'd63072;
			2465: outdata = 32'd63071;
			2466: outdata = 32'd63070;
			2467: outdata = 32'd63069;
			2468: outdata = 32'd63068;
			2469: outdata = 32'd63067;
			2470: outdata = 32'd63066;
			2471: outdata = 32'd63065;
			2472: outdata = 32'd63064;
			2473: outdata = 32'd63063;
			2474: outdata = 32'd63062;
			2475: outdata = 32'd63061;
			2476: outdata = 32'd63060;
			2477: outdata = 32'd63059;
			2478: outdata = 32'd63058;
			2479: outdata = 32'd63057;
			2480: outdata = 32'd63056;
			2481: outdata = 32'd63055;
			2482: outdata = 32'd63054;
			2483: outdata = 32'd63053;
			2484: outdata = 32'd63052;
			2485: outdata = 32'd63051;
			2486: outdata = 32'd63050;
			2487: outdata = 32'd63049;
			2488: outdata = 32'd63048;
			2489: outdata = 32'd63047;
			2490: outdata = 32'd63046;
			2491: outdata = 32'd63045;
			2492: outdata = 32'd63044;
			2493: outdata = 32'd63043;
			2494: outdata = 32'd63042;
			2495: outdata = 32'd63041;
			2496: outdata = 32'd63040;
			2497: outdata = 32'd63039;
			2498: outdata = 32'd63038;
			2499: outdata = 32'd63037;
			2500: outdata = 32'd63036;
			2501: outdata = 32'd63035;
			2502: outdata = 32'd63034;
			2503: outdata = 32'd63033;
			2504: outdata = 32'd63032;
			2505: outdata = 32'd63031;
			2506: outdata = 32'd63030;
			2507: outdata = 32'd63029;
			2508: outdata = 32'd63028;
			2509: outdata = 32'd63027;
			2510: outdata = 32'd63026;
			2511: outdata = 32'd63025;
			2512: outdata = 32'd63024;
			2513: outdata = 32'd63023;
			2514: outdata = 32'd63022;
			2515: outdata = 32'd63021;
			2516: outdata = 32'd63020;
			2517: outdata = 32'd63019;
			2518: outdata = 32'd63018;
			2519: outdata = 32'd63017;
			2520: outdata = 32'd63016;
			2521: outdata = 32'd63015;
			2522: outdata = 32'd63014;
			2523: outdata = 32'd63013;
			2524: outdata = 32'd63012;
			2525: outdata = 32'd63011;
			2526: outdata = 32'd63010;
			2527: outdata = 32'd63009;
			2528: outdata = 32'd63008;
			2529: outdata = 32'd63007;
			2530: outdata = 32'd63006;
			2531: outdata = 32'd63005;
			2532: outdata = 32'd63004;
			2533: outdata = 32'd63003;
			2534: outdata = 32'd63002;
			2535: outdata = 32'd63001;
			2536: outdata = 32'd63000;
			2537: outdata = 32'd62999;
			2538: outdata = 32'd62998;
			2539: outdata = 32'd62997;
			2540: outdata = 32'd62996;
			2541: outdata = 32'd62995;
			2542: outdata = 32'd62994;
			2543: outdata = 32'd62993;
			2544: outdata = 32'd62992;
			2545: outdata = 32'd62991;
			2546: outdata = 32'd62990;
			2547: outdata = 32'd62989;
			2548: outdata = 32'd62988;
			2549: outdata = 32'd62987;
			2550: outdata = 32'd62986;
			2551: outdata = 32'd62985;
			2552: outdata = 32'd62984;
			2553: outdata = 32'd62983;
			2554: outdata = 32'd62982;
			2555: outdata = 32'd62981;
			2556: outdata = 32'd62980;
			2557: outdata = 32'd62979;
			2558: outdata = 32'd62978;
			2559: outdata = 32'd62977;
			2560: outdata = 32'd62976;
			2561: outdata = 32'd62975;
			2562: outdata = 32'd62974;
			2563: outdata = 32'd62973;
			2564: outdata = 32'd62972;
			2565: outdata = 32'd62971;
			2566: outdata = 32'd62970;
			2567: outdata = 32'd62969;
			2568: outdata = 32'd62968;
			2569: outdata = 32'd62967;
			2570: outdata = 32'd62966;
			2571: outdata = 32'd62965;
			2572: outdata = 32'd62964;
			2573: outdata = 32'd62963;
			2574: outdata = 32'd62962;
			2575: outdata = 32'd62961;
			2576: outdata = 32'd62960;
			2577: outdata = 32'd62959;
			2578: outdata = 32'd62958;
			2579: outdata = 32'd62957;
			2580: outdata = 32'd62956;
			2581: outdata = 32'd62955;
			2582: outdata = 32'd62954;
			2583: outdata = 32'd62953;
			2584: outdata = 32'd62952;
			2585: outdata = 32'd62951;
			2586: outdata = 32'd62950;
			2587: outdata = 32'd62949;
			2588: outdata = 32'd62948;
			2589: outdata = 32'd62947;
			2590: outdata = 32'd62946;
			2591: outdata = 32'd62945;
			2592: outdata = 32'd62944;
			2593: outdata = 32'd62943;
			2594: outdata = 32'd62942;
			2595: outdata = 32'd62941;
			2596: outdata = 32'd62940;
			2597: outdata = 32'd62939;
			2598: outdata = 32'd62938;
			2599: outdata = 32'd62937;
			2600: outdata = 32'd62936;
			2601: outdata = 32'd62935;
			2602: outdata = 32'd62934;
			2603: outdata = 32'd62933;
			2604: outdata = 32'd62932;
			2605: outdata = 32'd62931;
			2606: outdata = 32'd62930;
			2607: outdata = 32'd62929;
			2608: outdata = 32'd62928;
			2609: outdata = 32'd62927;
			2610: outdata = 32'd62926;
			2611: outdata = 32'd62925;
			2612: outdata = 32'd62924;
			2613: outdata = 32'd62923;
			2614: outdata = 32'd62922;
			2615: outdata = 32'd62921;
			2616: outdata = 32'd62920;
			2617: outdata = 32'd62919;
			2618: outdata = 32'd62918;
			2619: outdata = 32'd62917;
			2620: outdata = 32'd62916;
			2621: outdata = 32'd62915;
			2622: outdata = 32'd62914;
			2623: outdata = 32'd62913;
			2624: outdata = 32'd62912;
			2625: outdata = 32'd62911;
			2626: outdata = 32'd62910;
			2627: outdata = 32'd62909;
			2628: outdata = 32'd62908;
			2629: outdata = 32'd62907;
			2630: outdata = 32'd62906;
			2631: outdata = 32'd62905;
			2632: outdata = 32'd62904;
			2633: outdata = 32'd62903;
			2634: outdata = 32'd62902;
			2635: outdata = 32'd62901;
			2636: outdata = 32'd62900;
			2637: outdata = 32'd62899;
			2638: outdata = 32'd62898;
			2639: outdata = 32'd62897;
			2640: outdata = 32'd62896;
			2641: outdata = 32'd62895;
			2642: outdata = 32'd62894;
			2643: outdata = 32'd62893;
			2644: outdata = 32'd62892;
			2645: outdata = 32'd62891;
			2646: outdata = 32'd62890;
			2647: outdata = 32'd62889;
			2648: outdata = 32'd62888;
			2649: outdata = 32'd62887;
			2650: outdata = 32'd62886;
			2651: outdata = 32'd62885;
			2652: outdata = 32'd62884;
			2653: outdata = 32'd62883;
			2654: outdata = 32'd62882;
			2655: outdata = 32'd62881;
			2656: outdata = 32'd62880;
			2657: outdata = 32'd62879;
			2658: outdata = 32'd62878;
			2659: outdata = 32'd62877;
			2660: outdata = 32'd62876;
			2661: outdata = 32'd62875;
			2662: outdata = 32'd62874;
			2663: outdata = 32'd62873;
			2664: outdata = 32'd62872;
			2665: outdata = 32'd62871;
			2666: outdata = 32'd62870;
			2667: outdata = 32'd62869;
			2668: outdata = 32'd62868;
			2669: outdata = 32'd62867;
			2670: outdata = 32'd62866;
			2671: outdata = 32'd62865;
			2672: outdata = 32'd62864;
			2673: outdata = 32'd62863;
			2674: outdata = 32'd62862;
			2675: outdata = 32'd62861;
			2676: outdata = 32'd62860;
			2677: outdata = 32'd62859;
			2678: outdata = 32'd62858;
			2679: outdata = 32'd62857;
			2680: outdata = 32'd62856;
			2681: outdata = 32'd62855;
			2682: outdata = 32'd62854;
			2683: outdata = 32'd62853;
			2684: outdata = 32'd62852;
			2685: outdata = 32'd62851;
			2686: outdata = 32'd62850;
			2687: outdata = 32'd62849;
			2688: outdata = 32'd62848;
			2689: outdata = 32'd62847;
			2690: outdata = 32'd62846;
			2691: outdata = 32'd62845;
			2692: outdata = 32'd62844;
			2693: outdata = 32'd62843;
			2694: outdata = 32'd62842;
			2695: outdata = 32'd62841;
			2696: outdata = 32'd62840;
			2697: outdata = 32'd62839;
			2698: outdata = 32'd62838;
			2699: outdata = 32'd62837;
			2700: outdata = 32'd62836;
			2701: outdata = 32'd62835;
			2702: outdata = 32'd62834;
			2703: outdata = 32'd62833;
			2704: outdata = 32'd62832;
			2705: outdata = 32'd62831;
			2706: outdata = 32'd62830;
			2707: outdata = 32'd62829;
			2708: outdata = 32'd62828;
			2709: outdata = 32'd62827;
			2710: outdata = 32'd62826;
			2711: outdata = 32'd62825;
			2712: outdata = 32'd62824;
			2713: outdata = 32'd62823;
			2714: outdata = 32'd62822;
			2715: outdata = 32'd62821;
			2716: outdata = 32'd62820;
			2717: outdata = 32'd62819;
			2718: outdata = 32'd62818;
			2719: outdata = 32'd62817;
			2720: outdata = 32'd62816;
			2721: outdata = 32'd62815;
			2722: outdata = 32'd62814;
			2723: outdata = 32'd62813;
			2724: outdata = 32'd62812;
			2725: outdata = 32'd62811;
			2726: outdata = 32'd62810;
			2727: outdata = 32'd62809;
			2728: outdata = 32'd62808;
			2729: outdata = 32'd62807;
			2730: outdata = 32'd62806;
			2731: outdata = 32'd62805;
			2732: outdata = 32'd62804;
			2733: outdata = 32'd62803;
			2734: outdata = 32'd62802;
			2735: outdata = 32'd62801;
			2736: outdata = 32'd62800;
			2737: outdata = 32'd62799;
			2738: outdata = 32'd62798;
			2739: outdata = 32'd62797;
			2740: outdata = 32'd62796;
			2741: outdata = 32'd62795;
			2742: outdata = 32'd62794;
			2743: outdata = 32'd62793;
			2744: outdata = 32'd62792;
			2745: outdata = 32'd62791;
			2746: outdata = 32'd62790;
			2747: outdata = 32'd62789;
			2748: outdata = 32'd62788;
			2749: outdata = 32'd62787;
			2750: outdata = 32'd62786;
			2751: outdata = 32'd62785;
			2752: outdata = 32'd62784;
			2753: outdata = 32'd62783;
			2754: outdata = 32'd62782;
			2755: outdata = 32'd62781;
			2756: outdata = 32'd62780;
			2757: outdata = 32'd62779;
			2758: outdata = 32'd62778;
			2759: outdata = 32'd62777;
			2760: outdata = 32'd62776;
			2761: outdata = 32'd62775;
			2762: outdata = 32'd62774;
			2763: outdata = 32'd62773;
			2764: outdata = 32'd62772;
			2765: outdata = 32'd62771;
			2766: outdata = 32'd62770;
			2767: outdata = 32'd62769;
			2768: outdata = 32'd62768;
			2769: outdata = 32'd62767;
			2770: outdata = 32'd62766;
			2771: outdata = 32'd62765;
			2772: outdata = 32'd62764;
			2773: outdata = 32'd62763;
			2774: outdata = 32'd62762;
			2775: outdata = 32'd62761;
			2776: outdata = 32'd62760;
			2777: outdata = 32'd62759;
			2778: outdata = 32'd62758;
			2779: outdata = 32'd62757;
			2780: outdata = 32'd62756;
			2781: outdata = 32'd62755;
			2782: outdata = 32'd62754;
			2783: outdata = 32'd62753;
			2784: outdata = 32'd62752;
			2785: outdata = 32'd62751;
			2786: outdata = 32'd62750;
			2787: outdata = 32'd62749;
			2788: outdata = 32'd62748;
			2789: outdata = 32'd62747;
			2790: outdata = 32'd62746;
			2791: outdata = 32'd62745;
			2792: outdata = 32'd62744;
			2793: outdata = 32'd62743;
			2794: outdata = 32'd62742;
			2795: outdata = 32'd62741;
			2796: outdata = 32'd62740;
			2797: outdata = 32'd62739;
			2798: outdata = 32'd62738;
			2799: outdata = 32'd62737;
			2800: outdata = 32'd62736;
			2801: outdata = 32'd62735;
			2802: outdata = 32'd62734;
			2803: outdata = 32'd62733;
			2804: outdata = 32'd62732;
			2805: outdata = 32'd62731;
			2806: outdata = 32'd62730;
			2807: outdata = 32'd62729;
			2808: outdata = 32'd62728;
			2809: outdata = 32'd62727;
			2810: outdata = 32'd62726;
			2811: outdata = 32'd62725;
			2812: outdata = 32'd62724;
			2813: outdata = 32'd62723;
			2814: outdata = 32'd62722;
			2815: outdata = 32'd62721;
			2816: outdata = 32'd62720;
			2817: outdata = 32'd62719;
			2818: outdata = 32'd62718;
			2819: outdata = 32'd62717;
			2820: outdata = 32'd62716;
			2821: outdata = 32'd62715;
			2822: outdata = 32'd62714;
			2823: outdata = 32'd62713;
			2824: outdata = 32'd62712;
			2825: outdata = 32'd62711;
			2826: outdata = 32'd62710;
			2827: outdata = 32'd62709;
			2828: outdata = 32'd62708;
			2829: outdata = 32'd62707;
			2830: outdata = 32'd62706;
			2831: outdata = 32'd62705;
			2832: outdata = 32'd62704;
			2833: outdata = 32'd62703;
			2834: outdata = 32'd62702;
			2835: outdata = 32'd62701;
			2836: outdata = 32'd62700;
			2837: outdata = 32'd62699;
			2838: outdata = 32'd62698;
			2839: outdata = 32'd62697;
			2840: outdata = 32'd62696;
			2841: outdata = 32'd62695;
			2842: outdata = 32'd62694;
			2843: outdata = 32'd62693;
			2844: outdata = 32'd62692;
			2845: outdata = 32'd62691;
			2846: outdata = 32'd62690;
			2847: outdata = 32'd62689;
			2848: outdata = 32'd62688;
			2849: outdata = 32'd62687;
			2850: outdata = 32'd62686;
			2851: outdata = 32'd62685;
			2852: outdata = 32'd62684;
			2853: outdata = 32'd62683;
			2854: outdata = 32'd62682;
			2855: outdata = 32'd62681;
			2856: outdata = 32'd62680;
			2857: outdata = 32'd62679;
			2858: outdata = 32'd62678;
			2859: outdata = 32'd62677;
			2860: outdata = 32'd62676;
			2861: outdata = 32'd62675;
			2862: outdata = 32'd62674;
			2863: outdata = 32'd62673;
			2864: outdata = 32'd62672;
			2865: outdata = 32'd62671;
			2866: outdata = 32'd62670;
			2867: outdata = 32'd62669;
			2868: outdata = 32'd62668;
			2869: outdata = 32'd62667;
			2870: outdata = 32'd62666;
			2871: outdata = 32'd62665;
			2872: outdata = 32'd62664;
			2873: outdata = 32'd62663;
			2874: outdata = 32'd62662;
			2875: outdata = 32'd62661;
			2876: outdata = 32'd62660;
			2877: outdata = 32'd62659;
			2878: outdata = 32'd62658;
			2879: outdata = 32'd62657;
			2880: outdata = 32'd62656;
			2881: outdata = 32'd62655;
			2882: outdata = 32'd62654;
			2883: outdata = 32'd62653;
			2884: outdata = 32'd62652;
			2885: outdata = 32'd62651;
			2886: outdata = 32'd62650;
			2887: outdata = 32'd62649;
			2888: outdata = 32'd62648;
			2889: outdata = 32'd62647;
			2890: outdata = 32'd62646;
			2891: outdata = 32'd62645;
			2892: outdata = 32'd62644;
			2893: outdata = 32'd62643;
			2894: outdata = 32'd62642;
			2895: outdata = 32'd62641;
			2896: outdata = 32'd62640;
			2897: outdata = 32'd62639;
			2898: outdata = 32'd62638;
			2899: outdata = 32'd62637;
			2900: outdata = 32'd62636;
			2901: outdata = 32'd62635;
			2902: outdata = 32'd62634;
			2903: outdata = 32'd62633;
			2904: outdata = 32'd62632;
			2905: outdata = 32'd62631;
			2906: outdata = 32'd62630;
			2907: outdata = 32'd62629;
			2908: outdata = 32'd62628;
			2909: outdata = 32'd62627;
			2910: outdata = 32'd62626;
			2911: outdata = 32'd62625;
			2912: outdata = 32'd62624;
			2913: outdata = 32'd62623;
			2914: outdata = 32'd62622;
			2915: outdata = 32'd62621;
			2916: outdata = 32'd62620;
			2917: outdata = 32'd62619;
			2918: outdata = 32'd62618;
			2919: outdata = 32'd62617;
			2920: outdata = 32'd62616;
			2921: outdata = 32'd62615;
			2922: outdata = 32'd62614;
			2923: outdata = 32'd62613;
			2924: outdata = 32'd62612;
			2925: outdata = 32'd62611;
			2926: outdata = 32'd62610;
			2927: outdata = 32'd62609;
			2928: outdata = 32'd62608;
			2929: outdata = 32'd62607;
			2930: outdata = 32'd62606;
			2931: outdata = 32'd62605;
			2932: outdata = 32'd62604;
			2933: outdata = 32'd62603;
			2934: outdata = 32'd62602;
			2935: outdata = 32'd62601;
			2936: outdata = 32'd62600;
			2937: outdata = 32'd62599;
			2938: outdata = 32'd62598;
			2939: outdata = 32'd62597;
			2940: outdata = 32'd62596;
			2941: outdata = 32'd62595;
			2942: outdata = 32'd62594;
			2943: outdata = 32'd62593;
			2944: outdata = 32'd62592;
			2945: outdata = 32'd62591;
			2946: outdata = 32'd62590;
			2947: outdata = 32'd62589;
			2948: outdata = 32'd62588;
			2949: outdata = 32'd62587;
			2950: outdata = 32'd62586;
			2951: outdata = 32'd62585;
			2952: outdata = 32'd62584;
			2953: outdata = 32'd62583;
			2954: outdata = 32'd62582;
			2955: outdata = 32'd62581;
			2956: outdata = 32'd62580;
			2957: outdata = 32'd62579;
			2958: outdata = 32'd62578;
			2959: outdata = 32'd62577;
			2960: outdata = 32'd62576;
			2961: outdata = 32'd62575;
			2962: outdata = 32'd62574;
			2963: outdata = 32'd62573;
			2964: outdata = 32'd62572;
			2965: outdata = 32'd62571;
			2966: outdata = 32'd62570;
			2967: outdata = 32'd62569;
			2968: outdata = 32'd62568;
			2969: outdata = 32'd62567;
			2970: outdata = 32'd62566;
			2971: outdata = 32'd62565;
			2972: outdata = 32'd62564;
			2973: outdata = 32'd62563;
			2974: outdata = 32'd62562;
			2975: outdata = 32'd62561;
			2976: outdata = 32'd62560;
			2977: outdata = 32'd62559;
			2978: outdata = 32'd62558;
			2979: outdata = 32'd62557;
			2980: outdata = 32'd62556;
			2981: outdata = 32'd62555;
			2982: outdata = 32'd62554;
			2983: outdata = 32'd62553;
			2984: outdata = 32'd62552;
			2985: outdata = 32'd62551;
			2986: outdata = 32'd62550;
			2987: outdata = 32'd62549;
			2988: outdata = 32'd62548;
			2989: outdata = 32'd62547;
			2990: outdata = 32'd62546;
			2991: outdata = 32'd62545;
			2992: outdata = 32'd62544;
			2993: outdata = 32'd62543;
			2994: outdata = 32'd62542;
			2995: outdata = 32'd62541;
			2996: outdata = 32'd62540;
			2997: outdata = 32'd62539;
			2998: outdata = 32'd62538;
			2999: outdata = 32'd62537;
			3000: outdata = 32'd62536;
			3001: outdata = 32'd62535;
			3002: outdata = 32'd62534;
			3003: outdata = 32'd62533;
			3004: outdata = 32'd62532;
			3005: outdata = 32'd62531;
			3006: outdata = 32'd62530;
			3007: outdata = 32'd62529;
			3008: outdata = 32'd62528;
			3009: outdata = 32'd62527;
			3010: outdata = 32'd62526;
			3011: outdata = 32'd62525;
			3012: outdata = 32'd62524;
			3013: outdata = 32'd62523;
			3014: outdata = 32'd62522;
			3015: outdata = 32'd62521;
			3016: outdata = 32'd62520;
			3017: outdata = 32'd62519;
			3018: outdata = 32'd62518;
			3019: outdata = 32'd62517;
			3020: outdata = 32'd62516;
			3021: outdata = 32'd62515;
			3022: outdata = 32'd62514;
			3023: outdata = 32'd62513;
			3024: outdata = 32'd62512;
			3025: outdata = 32'd62511;
			3026: outdata = 32'd62510;
			3027: outdata = 32'd62509;
			3028: outdata = 32'd62508;
			3029: outdata = 32'd62507;
			3030: outdata = 32'd62506;
			3031: outdata = 32'd62505;
			3032: outdata = 32'd62504;
			3033: outdata = 32'd62503;
			3034: outdata = 32'd62502;
			3035: outdata = 32'd62501;
			3036: outdata = 32'd62500;
			3037: outdata = 32'd62499;
			3038: outdata = 32'd62498;
			3039: outdata = 32'd62497;
			3040: outdata = 32'd62496;
			3041: outdata = 32'd62495;
			3042: outdata = 32'd62494;
			3043: outdata = 32'd62493;
			3044: outdata = 32'd62492;
			3045: outdata = 32'd62491;
			3046: outdata = 32'd62490;
			3047: outdata = 32'd62489;
			3048: outdata = 32'd62488;
			3049: outdata = 32'd62487;
			3050: outdata = 32'd62486;
			3051: outdata = 32'd62485;
			3052: outdata = 32'd62484;
			3053: outdata = 32'd62483;
			3054: outdata = 32'd62482;
			3055: outdata = 32'd62481;
			3056: outdata = 32'd62480;
			3057: outdata = 32'd62479;
			3058: outdata = 32'd62478;
			3059: outdata = 32'd62477;
			3060: outdata = 32'd62476;
			3061: outdata = 32'd62475;
			3062: outdata = 32'd62474;
			3063: outdata = 32'd62473;
			3064: outdata = 32'd62472;
			3065: outdata = 32'd62471;
			3066: outdata = 32'd62470;
			3067: outdata = 32'd62469;
			3068: outdata = 32'd62468;
			3069: outdata = 32'd62467;
			3070: outdata = 32'd62466;
			3071: outdata = 32'd62465;
			3072: outdata = 32'd62464;
			3073: outdata = 32'd62463;
			3074: outdata = 32'd62462;
			3075: outdata = 32'd62461;
			3076: outdata = 32'd62460;
			3077: outdata = 32'd62459;
			3078: outdata = 32'd62458;
			3079: outdata = 32'd62457;
			3080: outdata = 32'd62456;
			3081: outdata = 32'd62455;
			3082: outdata = 32'd62454;
			3083: outdata = 32'd62453;
			3084: outdata = 32'd62452;
			3085: outdata = 32'd62451;
			3086: outdata = 32'd62450;
			3087: outdata = 32'd62449;
			3088: outdata = 32'd62448;
			3089: outdata = 32'd62447;
			3090: outdata = 32'd62446;
			3091: outdata = 32'd62445;
			3092: outdata = 32'd62444;
			3093: outdata = 32'd62443;
			3094: outdata = 32'd62442;
			3095: outdata = 32'd62441;
			3096: outdata = 32'd62440;
			3097: outdata = 32'd62439;
			3098: outdata = 32'd62438;
			3099: outdata = 32'd62437;
			3100: outdata = 32'd62436;
			3101: outdata = 32'd62435;
			3102: outdata = 32'd62434;
			3103: outdata = 32'd62433;
			3104: outdata = 32'd62432;
			3105: outdata = 32'd62431;
			3106: outdata = 32'd62430;
			3107: outdata = 32'd62429;
			3108: outdata = 32'd62428;
			3109: outdata = 32'd62427;
			3110: outdata = 32'd62426;
			3111: outdata = 32'd62425;
			3112: outdata = 32'd62424;
			3113: outdata = 32'd62423;
			3114: outdata = 32'd62422;
			3115: outdata = 32'd62421;
			3116: outdata = 32'd62420;
			3117: outdata = 32'd62419;
			3118: outdata = 32'd62418;
			3119: outdata = 32'd62417;
			3120: outdata = 32'd62416;
			3121: outdata = 32'd62415;
			3122: outdata = 32'd62414;
			3123: outdata = 32'd62413;
			3124: outdata = 32'd62412;
			3125: outdata = 32'd62411;
			3126: outdata = 32'd62410;
			3127: outdata = 32'd62409;
			3128: outdata = 32'd62408;
			3129: outdata = 32'd62407;
			3130: outdata = 32'd62406;
			3131: outdata = 32'd62405;
			3132: outdata = 32'd62404;
			3133: outdata = 32'd62403;
			3134: outdata = 32'd62402;
			3135: outdata = 32'd62401;
			3136: outdata = 32'd62400;
			3137: outdata = 32'd62399;
			3138: outdata = 32'd62398;
			3139: outdata = 32'd62397;
			3140: outdata = 32'd62396;
			3141: outdata = 32'd62395;
			3142: outdata = 32'd62394;
			3143: outdata = 32'd62393;
			3144: outdata = 32'd62392;
			3145: outdata = 32'd62391;
			3146: outdata = 32'd62390;
			3147: outdata = 32'd62389;
			3148: outdata = 32'd62388;
			3149: outdata = 32'd62387;
			3150: outdata = 32'd62386;
			3151: outdata = 32'd62385;
			3152: outdata = 32'd62384;
			3153: outdata = 32'd62383;
			3154: outdata = 32'd62382;
			3155: outdata = 32'd62381;
			3156: outdata = 32'd62380;
			3157: outdata = 32'd62379;
			3158: outdata = 32'd62378;
			3159: outdata = 32'd62377;
			3160: outdata = 32'd62376;
			3161: outdata = 32'd62375;
			3162: outdata = 32'd62374;
			3163: outdata = 32'd62373;
			3164: outdata = 32'd62372;
			3165: outdata = 32'd62371;
			3166: outdata = 32'd62370;
			3167: outdata = 32'd62369;
			3168: outdata = 32'd62368;
			3169: outdata = 32'd62367;
			3170: outdata = 32'd62366;
			3171: outdata = 32'd62365;
			3172: outdata = 32'd62364;
			3173: outdata = 32'd62363;
			3174: outdata = 32'd62362;
			3175: outdata = 32'd62361;
			3176: outdata = 32'd62360;
			3177: outdata = 32'd62359;
			3178: outdata = 32'd62358;
			3179: outdata = 32'd62357;
			3180: outdata = 32'd62356;
			3181: outdata = 32'd62355;
			3182: outdata = 32'd62354;
			3183: outdata = 32'd62353;
			3184: outdata = 32'd62352;
			3185: outdata = 32'd62351;
			3186: outdata = 32'd62350;
			3187: outdata = 32'd62349;
			3188: outdata = 32'd62348;
			3189: outdata = 32'd62347;
			3190: outdata = 32'd62346;
			3191: outdata = 32'd62345;
			3192: outdata = 32'd62344;
			3193: outdata = 32'd62343;
			3194: outdata = 32'd62342;
			3195: outdata = 32'd62341;
			3196: outdata = 32'd62340;
			3197: outdata = 32'd62339;
			3198: outdata = 32'd62338;
			3199: outdata = 32'd62337;
			3200: outdata = 32'd62336;
			3201: outdata = 32'd62335;
			3202: outdata = 32'd62334;
			3203: outdata = 32'd62333;
			3204: outdata = 32'd62332;
			3205: outdata = 32'd62331;
			3206: outdata = 32'd62330;
			3207: outdata = 32'd62329;
			3208: outdata = 32'd62328;
			3209: outdata = 32'd62327;
			3210: outdata = 32'd62326;
			3211: outdata = 32'd62325;
			3212: outdata = 32'd62324;
			3213: outdata = 32'd62323;
			3214: outdata = 32'd62322;
			3215: outdata = 32'd62321;
			3216: outdata = 32'd62320;
			3217: outdata = 32'd62319;
			3218: outdata = 32'd62318;
			3219: outdata = 32'd62317;
			3220: outdata = 32'd62316;
			3221: outdata = 32'd62315;
			3222: outdata = 32'd62314;
			3223: outdata = 32'd62313;
			3224: outdata = 32'd62312;
			3225: outdata = 32'd62311;
			3226: outdata = 32'd62310;
			3227: outdata = 32'd62309;
			3228: outdata = 32'd62308;
			3229: outdata = 32'd62307;
			3230: outdata = 32'd62306;
			3231: outdata = 32'd62305;
			3232: outdata = 32'd62304;
			3233: outdata = 32'd62303;
			3234: outdata = 32'd62302;
			3235: outdata = 32'd62301;
			3236: outdata = 32'd62300;
			3237: outdata = 32'd62299;
			3238: outdata = 32'd62298;
			3239: outdata = 32'd62297;
			3240: outdata = 32'd62296;
			3241: outdata = 32'd62295;
			3242: outdata = 32'd62294;
			3243: outdata = 32'd62293;
			3244: outdata = 32'd62292;
			3245: outdata = 32'd62291;
			3246: outdata = 32'd62290;
			3247: outdata = 32'd62289;
			3248: outdata = 32'd62288;
			3249: outdata = 32'd62287;
			3250: outdata = 32'd62286;
			3251: outdata = 32'd62285;
			3252: outdata = 32'd62284;
			3253: outdata = 32'd62283;
			3254: outdata = 32'd62282;
			3255: outdata = 32'd62281;
			3256: outdata = 32'd62280;
			3257: outdata = 32'd62279;
			3258: outdata = 32'd62278;
			3259: outdata = 32'd62277;
			3260: outdata = 32'd62276;
			3261: outdata = 32'd62275;
			3262: outdata = 32'd62274;
			3263: outdata = 32'd62273;
			3264: outdata = 32'd62272;
			3265: outdata = 32'd62271;
			3266: outdata = 32'd62270;
			3267: outdata = 32'd62269;
			3268: outdata = 32'd62268;
			3269: outdata = 32'd62267;
			3270: outdata = 32'd62266;
			3271: outdata = 32'd62265;
			3272: outdata = 32'd62264;
			3273: outdata = 32'd62263;
			3274: outdata = 32'd62262;
			3275: outdata = 32'd62261;
			3276: outdata = 32'd62260;
			3277: outdata = 32'd62259;
			3278: outdata = 32'd62258;
			3279: outdata = 32'd62257;
			3280: outdata = 32'd62256;
			3281: outdata = 32'd62255;
			3282: outdata = 32'd62254;
			3283: outdata = 32'd62253;
			3284: outdata = 32'd62252;
			3285: outdata = 32'd62251;
			3286: outdata = 32'd62250;
			3287: outdata = 32'd62249;
			3288: outdata = 32'd62248;
			3289: outdata = 32'd62247;
			3290: outdata = 32'd62246;
			3291: outdata = 32'd62245;
			3292: outdata = 32'd62244;
			3293: outdata = 32'd62243;
			3294: outdata = 32'd62242;
			3295: outdata = 32'd62241;
			3296: outdata = 32'd62240;
			3297: outdata = 32'd62239;
			3298: outdata = 32'd62238;
			3299: outdata = 32'd62237;
			3300: outdata = 32'd62236;
			3301: outdata = 32'd62235;
			3302: outdata = 32'd62234;
			3303: outdata = 32'd62233;
			3304: outdata = 32'd62232;
			3305: outdata = 32'd62231;
			3306: outdata = 32'd62230;
			3307: outdata = 32'd62229;
			3308: outdata = 32'd62228;
			3309: outdata = 32'd62227;
			3310: outdata = 32'd62226;
			3311: outdata = 32'd62225;
			3312: outdata = 32'd62224;
			3313: outdata = 32'd62223;
			3314: outdata = 32'd62222;
			3315: outdata = 32'd62221;
			3316: outdata = 32'd62220;
			3317: outdata = 32'd62219;
			3318: outdata = 32'd62218;
			3319: outdata = 32'd62217;
			3320: outdata = 32'd62216;
			3321: outdata = 32'd62215;
			3322: outdata = 32'd62214;
			3323: outdata = 32'd62213;
			3324: outdata = 32'd62212;
			3325: outdata = 32'd62211;
			3326: outdata = 32'd62210;
			3327: outdata = 32'd62209;
			3328: outdata = 32'd62208;
			3329: outdata = 32'd62207;
			3330: outdata = 32'd62206;
			3331: outdata = 32'd62205;
			3332: outdata = 32'd62204;
			3333: outdata = 32'd62203;
			3334: outdata = 32'd62202;
			3335: outdata = 32'd62201;
			3336: outdata = 32'd62200;
			3337: outdata = 32'd62199;
			3338: outdata = 32'd62198;
			3339: outdata = 32'd62197;
			3340: outdata = 32'd62196;
			3341: outdata = 32'd62195;
			3342: outdata = 32'd62194;
			3343: outdata = 32'd62193;
			3344: outdata = 32'd62192;
			3345: outdata = 32'd62191;
			3346: outdata = 32'd62190;
			3347: outdata = 32'd62189;
			3348: outdata = 32'd62188;
			3349: outdata = 32'd62187;
			3350: outdata = 32'd62186;
			3351: outdata = 32'd62185;
			3352: outdata = 32'd62184;
			3353: outdata = 32'd62183;
			3354: outdata = 32'd62182;
			3355: outdata = 32'd62181;
			3356: outdata = 32'd62180;
			3357: outdata = 32'd62179;
			3358: outdata = 32'd62178;
			3359: outdata = 32'd62177;
			3360: outdata = 32'd62176;
			3361: outdata = 32'd62175;
			3362: outdata = 32'd62174;
			3363: outdata = 32'd62173;
			3364: outdata = 32'd62172;
			3365: outdata = 32'd62171;
			3366: outdata = 32'd62170;
			3367: outdata = 32'd62169;
			3368: outdata = 32'd62168;
			3369: outdata = 32'd62167;
			3370: outdata = 32'd62166;
			3371: outdata = 32'd62165;
			3372: outdata = 32'd62164;
			3373: outdata = 32'd62163;
			3374: outdata = 32'd62162;
			3375: outdata = 32'd62161;
			3376: outdata = 32'd62160;
			3377: outdata = 32'd62159;
			3378: outdata = 32'd62158;
			3379: outdata = 32'd62157;
			3380: outdata = 32'd62156;
			3381: outdata = 32'd62155;
			3382: outdata = 32'd62154;
			3383: outdata = 32'd62153;
			3384: outdata = 32'd62152;
			3385: outdata = 32'd62151;
			3386: outdata = 32'd62150;
			3387: outdata = 32'd62149;
			3388: outdata = 32'd62148;
			3389: outdata = 32'd62147;
			3390: outdata = 32'd62146;
			3391: outdata = 32'd62145;
			3392: outdata = 32'd62144;
			3393: outdata = 32'd62143;
			3394: outdata = 32'd62142;
			3395: outdata = 32'd62141;
			3396: outdata = 32'd62140;
			3397: outdata = 32'd62139;
			3398: outdata = 32'd62138;
			3399: outdata = 32'd62137;
			3400: outdata = 32'd62136;
			3401: outdata = 32'd62135;
			3402: outdata = 32'd62134;
			3403: outdata = 32'd62133;
			3404: outdata = 32'd62132;
			3405: outdata = 32'd62131;
			3406: outdata = 32'd62130;
			3407: outdata = 32'd62129;
			3408: outdata = 32'd62128;
			3409: outdata = 32'd62127;
			3410: outdata = 32'd62126;
			3411: outdata = 32'd62125;
			3412: outdata = 32'd62124;
			3413: outdata = 32'd62123;
			3414: outdata = 32'd62122;
			3415: outdata = 32'd62121;
			3416: outdata = 32'd62120;
			3417: outdata = 32'd62119;
			3418: outdata = 32'd62118;
			3419: outdata = 32'd62117;
			3420: outdata = 32'd62116;
			3421: outdata = 32'd62115;
			3422: outdata = 32'd62114;
			3423: outdata = 32'd62113;
			3424: outdata = 32'd62112;
			3425: outdata = 32'd62111;
			3426: outdata = 32'd62110;
			3427: outdata = 32'd62109;
			3428: outdata = 32'd62108;
			3429: outdata = 32'd62107;
			3430: outdata = 32'd62106;
			3431: outdata = 32'd62105;
			3432: outdata = 32'd62104;
			3433: outdata = 32'd62103;
			3434: outdata = 32'd62102;
			3435: outdata = 32'd62101;
			3436: outdata = 32'd62100;
			3437: outdata = 32'd62099;
			3438: outdata = 32'd62098;
			3439: outdata = 32'd62097;
			3440: outdata = 32'd62096;
			3441: outdata = 32'd62095;
			3442: outdata = 32'd62094;
			3443: outdata = 32'd62093;
			3444: outdata = 32'd62092;
			3445: outdata = 32'd62091;
			3446: outdata = 32'd62090;
			3447: outdata = 32'd62089;
			3448: outdata = 32'd62088;
			3449: outdata = 32'd62087;
			3450: outdata = 32'd62086;
			3451: outdata = 32'd62085;
			3452: outdata = 32'd62084;
			3453: outdata = 32'd62083;
			3454: outdata = 32'd62082;
			3455: outdata = 32'd62081;
			3456: outdata = 32'd62080;
			3457: outdata = 32'd62079;
			3458: outdata = 32'd62078;
			3459: outdata = 32'd62077;
			3460: outdata = 32'd62076;
			3461: outdata = 32'd62075;
			3462: outdata = 32'd62074;
			3463: outdata = 32'd62073;
			3464: outdata = 32'd62072;
			3465: outdata = 32'd62071;
			3466: outdata = 32'd62070;
			3467: outdata = 32'd62069;
			3468: outdata = 32'd62068;
			3469: outdata = 32'd62067;
			3470: outdata = 32'd62066;
			3471: outdata = 32'd62065;
			3472: outdata = 32'd62064;
			3473: outdata = 32'd62063;
			3474: outdata = 32'd62062;
			3475: outdata = 32'd62061;
			3476: outdata = 32'd62060;
			3477: outdata = 32'd62059;
			3478: outdata = 32'd62058;
			3479: outdata = 32'd62057;
			3480: outdata = 32'd62056;
			3481: outdata = 32'd62055;
			3482: outdata = 32'd62054;
			3483: outdata = 32'd62053;
			3484: outdata = 32'd62052;
			3485: outdata = 32'd62051;
			3486: outdata = 32'd62050;
			3487: outdata = 32'd62049;
			3488: outdata = 32'd62048;
			3489: outdata = 32'd62047;
			3490: outdata = 32'd62046;
			3491: outdata = 32'd62045;
			3492: outdata = 32'd62044;
			3493: outdata = 32'd62043;
			3494: outdata = 32'd62042;
			3495: outdata = 32'd62041;
			3496: outdata = 32'd62040;
			3497: outdata = 32'd62039;
			3498: outdata = 32'd62038;
			3499: outdata = 32'd62037;
			3500: outdata = 32'd62036;
			3501: outdata = 32'd62035;
			3502: outdata = 32'd62034;
			3503: outdata = 32'd62033;
			3504: outdata = 32'd62032;
			3505: outdata = 32'd62031;
			3506: outdata = 32'd62030;
			3507: outdata = 32'd62029;
			3508: outdata = 32'd62028;
			3509: outdata = 32'd62027;
			3510: outdata = 32'd62026;
			3511: outdata = 32'd62025;
			3512: outdata = 32'd62024;
			3513: outdata = 32'd62023;
			3514: outdata = 32'd62022;
			3515: outdata = 32'd62021;
			3516: outdata = 32'd62020;
			3517: outdata = 32'd62019;
			3518: outdata = 32'd62018;
			3519: outdata = 32'd62017;
			3520: outdata = 32'd62016;
			3521: outdata = 32'd62015;
			3522: outdata = 32'd62014;
			3523: outdata = 32'd62013;
			3524: outdata = 32'd62012;
			3525: outdata = 32'd62011;
			3526: outdata = 32'd62010;
			3527: outdata = 32'd62009;
			3528: outdata = 32'd62008;
			3529: outdata = 32'd62007;
			3530: outdata = 32'd62006;
			3531: outdata = 32'd62005;
			3532: outdata = 32'd62004;
			3533: outdata = 32'd62003;
			3534: outdata = 32'd62002;
			3535: outdata = 32'd62001;
			3536: outdata = 32'd62000;
			3537: outdata = 32'd61999;
			3538: outdata = 32'd61998;
			3539: outdata = 32'd61997;
			3540: outdata = 32'd61996;
			3541: outdata = 32'd61995;
			3542: outdata = 32'd61994;
			3543: outdata = 32'd61993;
			3544: outdata = 32'd61992;
			3545: outdata = 32'd61991;
			3546: outdata = 32'd61990;
			3547: outdata = 32'd61989;
			3548: outdata = 32'd61988;
			3549: outdata = 32'd61987;
			3550: outdata = 32'd61986;
			3551: outdata = 32'd61985;
			3552: outdata = 32'd61984;
			3553: outdata = 32'd61983;
			3554: outdata = 32'd61982;
			3555: outdata = 32'd61981;
			3556: outdata = 32'd61980;
			3557: outdata = 32'd61979;
			3558: outdata = 32'd61978;
			3559: outdata = 32'd61977;
			3560: outdata = 32'd61976;
			3561: outdata = 32'd61975;
			3562: outdata = 32'd61974;
			3563: outdata = 32'd61973;
			3564: outdata = 32'd61972;
			3565: outdata = 32'd61971;
			3566: outdata = 32'd61970;
			3567: outdata = 32'd61969;
			3568: outdata = 32'd61968;
			3569: outdata = 32'd61967;
			3570: outdata = 32'd61966;
			3571: outdata = 32'd61965;
			3572: outdata = 32'd61964;
			3573: outdata = 32'd61963;
			3574: outdata = 32'd61962;
			3575: outdata = 32'd61961;
			3576: outdata = 32'd61960;
			3577: outdata = 32'd61959;
			3578: outdata = 32'd61958;
			3579: outdata = 32'd61957;
			3580: outdata = 32'd61956;
			3581: outdata = 32'd61955;
			3582: outdata = 32'd61954;
			3583: outdata = 32'd61953;
			3584: outdata = 32'd61952;
			3585: outdata = 32'd61951;
			3586: outdata = 32'd61950;
			3587: outdata = 32'd61949;
			3588: outdata = 32'd61948;
			3589: outdata = 32'd61947;
			3590: outdata = 32'd61946;
			3591: outdata = 32'd61945;
			3592: outdata = 32'd61944;
			3593: outdata = 32'd61943;
			3594: outdata = 32'd61942;
			3595: outdata = 32'd61941;
			3596: outdata = 32'd61940;
			3597: outdata = 32'd61939;
			3598: outdata = 32'd61938;
			3599: outdata = 32'd61937;
			3600: outdata = 32'd61936;
			3601: outdata = 32'd61935;
			3602: outdata = 32'd61934;
			3603: outdata = 32'd61933;
			3604: outdata = 32'd61932;
			3605: outdata = 32'd61931;
			3606: outdata = 32'd61930;
			3607: outdata = 32'd61929;
			3608: outdata = 32'd61928;
			3609: outdata = 32'd61927;
			3610: outdata = 32'd61926;
			3611: outdata = 32'd61925;
			3612: outdata = 32'd61924;
			3613: outdata = 32'd61923;
			3614: outdata = 32'd61922;
			3615: outdata = 32'd61921;
			3616: outdata = 32'd61920;
			3617: outdata = 32'd61919;
			3618: outdata = 32'd61918;
			3619: outdata = 32'd61917;
			3620: outdata = 32'd61916;
			3621: outdata = 32'd61915;
			3622: outdata = 32'd61914;
			3623: outdata = 32'd61913;
			3624: outdata = 32'd61912;
			3625: outdata = 32'd61911;
			3626: outdata = 32'd61910;
			3627: outdata = 32'd61909;
			3628: outdata = 32'd61908;
			3629: outdata = 32'd61907;
			3630: outdata = 32'd61906;
			3631: outdata = 32'd61905;
			3632: outdata = 32'd61904;
			3633: outdata = 32'd61903;
			3634: outdata = 32'd61902;
			3635: outdata = 32'd61901;
			3636: outdata = 32'd61900;
			3637: outdata = 32'd61899;
			3638: outdata = 32'd61898;
			3639: outdata = 32'd61897;
			3640: outdata = 32'd61896;
			3641: outdata = 32'd61895;
			3642: outdata = 32'd61894;
			3643: outdata = 32'd61893;
			3644: outdata = 32'd61892;
			3645: outdata = 32'd61891;
			3646: outdata = 32'd61890;
			3647: outdata = 32'd61889;
			3648: outdata = 32'd61888;
			3649: outdata = 32'd61887;
			3650: outdata = 32'd61886;
			3651: outdata = 32'd61885;
			3652: outdata = 32'd61884;
			3653: outdata = 32'd61883;
			3654: outdata = 32'd61882;
			3655: outdata = 32'd61881;
			3656: outdata = 32'd61880;
			3657: outdata = 32'd61879;
			3658: outdata = 32'd61878;
			3659: outdata = 32'd61877;
			3660: outdata = 32'd61876;
			3661: outdata = 32'd61875;
			3662: outdata = 32'd61874;
			3663: outdata = 32'd61873;
			3664: outdata = 32'd61872;
			3665: outdata = 32'd61871;
			3666: outdata = 32'd61870;
			3667: outdata = 32'd61869;
			3668: outdata = 32'd61868;
			3669: outdata = 32'd61867;
			3670: outdata = 32'd61866;
			3671: outdata = 32'd61865;
			3672: outdata = 32'd61864;
			3673: outdata = 32'd61863;
			3674: outdata = 32'd61862;
			3675: outdata = 32'd61861;
			3676: outdata = 32'd61860;
			3677: outdata = 32'd61859;
			3678: outdata = 32'd61858;
			3679: outdata = 32'd61857;
			3680: outdata = 32'd61856;
			3681: outdata = 32'd61855;
			3682: outdata = 32'd61854;
			3683: outdata = 32'd61853;
			3684: outdata = 32'd61852;
			3685: outdata = 32'd61851;
			3686: outdata = 32'd61850;
			3687: outdata = 32'd61849;
			3688: outdata = 32'd61848;
			3689: outdata = 32'd61847;
			3690: outdata = 32'd61846;
			3691: outdata = 32'd61845;
			3692: outdata = 32'd61844;
			3693: outdata = 32'd61843;
			3694: outdata = 32'd61842;
			3695: outdata = 32'd61841;
			3696: outdata = 32'd61840;
			3697: outdata = 32'd61839;
			3698: outdata = 32'd61838;
			3699: outdata = 32'd61837;
			3700: outdata = 32'd61836;
			3701: outdata = 32'd61835;
			3702: outdata = 32'd61834;
			3703: outdata = 32'd61833;
			3704: outdata = 32'd61832;
			3705: outdata = 32'd61831;
			3706: outdata = 32'd61830;
			3707: outdata = 32'd61829;
			3708: outdata = 32'd61828;
			3709: outdata = 32'd61827;
			3710: outdata = 32'd61826;
			3711: outdata = 32'd61825;
			3712: outdata = 32'd61824;
			3713: outdata = 32'd61823;
			3714: outdata = 32'd61822;
			3715: outdata = 32'd61821;
			3716: outdata = 32'd61820;
			3717: outdata = 32'd61819;
			3718: outdata = 32'd61818;
			3719: outdata = 32'd61817;
			3720: outdata = 32'd61816;
			3721: outdata = 32'd61815;
			3722: outdata = 32'd61814;
			3723: outdata = 32'd61813;
			3724: outdata = 32'd61812;
			3725: outdata = 32'd61811;
			3726: outdata = 32'd61810;
			3727: outdata = 32'd61809;
			3728: outdata = 32'd61808;
			3729: outdata = 32'd61807;
			3730: outdata = 32'd61806;
			3731: outdata = 32'd61805;
			3732: outdata = 32'd61804;
			3733: outdata = 32'd61803;
			3734: outdata = 32'd61802;
			3735: outdata = 32'd61801;
			3736: outdata = 32'd61800;
			3737: outdata = 32'd61799;
			3738: outdata = 32'd61798;
			3739: outdata = 32'd61797;
			3740: outdata = 32'd61796;
			3741: outdata = 32'd61795;
			3742: outdata = 32'd61794;
			3743: outdata = 32'd61793;
			3744: outdata = 32'd61792;
			3745: outdata = 32'd61791;
			3746: outdata = 32'd61790;
			3747: outdata = 32'd61789;
			3748: outdata = 32'd61788;
			3749: outdata = 32'd61787;
			3750: outdata = 32'd61786;
			3751: outdata = 32'd61785;
			3752: outdata = 32'd61784;
			3753: outdata = 32'd61783;
			3754: outdata = 32'd61782;
			3755: outdata = 32'd61781;
			3756: outdata = 32'd61780;
			3757: outdata = 32'd61779;
			3758: outdata = 32'd61778;
			3759: outdata = 32'd61777;
			3760: outdata = 32'd61776;
			3761: outdata = 32'd61775;
			3762: outdata = 32'd61774;
			3763: outdata = 32'd61773;
			3764: outdata = 32'd61772;
			3765: outdata = 32'd61771;
			3766: outdata = 32'd61770;
			3767: outdata = 32'd61769;
			3768: outdata = 32'd61768;
			3769: outdata = 32'd61767;
			3770: outdata = 32'd61766;
			3771: outdata = 32'd61765;
			3772: outdata = 32'd61764;
			3773: outdata = 32'd61763;
			3774: outdata = 32'd61762;
			3775: outdata = 32'd61761;
			3776: outdata = 32'd61760;
			3777: outdata = 32'd61759;
			3778: outdata = 32'd61758;
			3779: outdata = 32'd61757;
			3780: outdata = 32'd61756;
			3781: outdata = 32'd61755;
			3782: outdata = 32'd61754;
			3783: outdata = 32'd61753;
			3784: outdata = 32'd61752;
			3785: outdata = 32'd61751;
			3786: outdata = 32'd61750;
			3787: outdata = 32'd61749;
			3788: outdata = 32'd61748;
			3789: outdata = 32'd61747;
			3790: outdata = 32'd61746;
			3791: outdata = 32'd61745;
			3792: outdata = 32'd61744;
			3793: outdata = 32'd61743;
			3794: outdata = 32'd61742;
			3795: outdata = 32'd61741;
			3796: outdata = 32'd61740;
			3797: outdata = 32'd61739;
			3798: outdata = 32'd61738;
			3799: outdata = 32'd61737;
			3800: outdata = 32'd61736;
			3801: outdata = 32'd61735;
			3802: outdata = 32'd61734;
			3803: outdata = 32'd61733;
			3804: outdata = 32'd61732;
			3805: outdata = 32'd61731;
			3806: outdata = 32'd61730;
			3807: outdata = 32'd61729;
			3808: outdata = 32'd61728;
			3809: outdata = 32'd61727;
			3810: outdata = 32'd61726;
			3811: outdata = 32'd61725;
			3812: outdata = 32'd61724;
			3813: outdata = 32'd61723;
			3814: outdata = 32'd61722;
			3815: outdata = 32'd61721;
			3816: outdata = 32'd61720;
			3817: outdata = 32'd61719;
			3818: outdata = 32'd61718;
			3819: outdata = 32'd61717;
			3820: outdata = 32'd61716;
			3821: outdata = 32'd61715;
			3822: outdata = 32'd61714;
			3823: outdata = 32'd61713;
			3824: outdata = 32'd61712;
			3825: outdata = 32'd61711;
			3826: outdata = 32'd61710;
			3827: outdata = 32'd61709;
			3828: outdata = 32'd61708;
			3829: outdata = 32'd61707;
			3830: outdata = 32'd61706;
			3831: outdata = 32'd61705;
			3832: outdata = 32'd61704;
			3833: outdata = 32'd61703;
			3834: outdata = 32'd61702;
			3835: outdata = 32'd61701;
			3836: outdata = 32'd61700;
			3837: outdata = 32'd61699;
			3838: outdata = 32'd61698;
			3839: outdata = 32'd61697;
			3840: outdata = 32'd61696;
			3841: outdata = 32'd61695;
			3842: outdata = 32'd61694;
			3843: outdata = 32'd61693;
			3844: outdata = 32'd61692;
			3845: outdata = 32'd61691;
			3846: outdata = 32'd61690;
			3847: outdata = 32'd61689;
			3848: outdata = 32'd61688;
			3849: outdata = 32'd61687;
			3850: outdata = 32'd61686;
			3851: outdata = 32'd61685;
			3852: outdata = 32'd61684;
			3853: outdata = 32'd61683;
			3854: outdata = 32'd61682;
			3855: outdata = 32'd61681;
			3856: outdata = 32'd61680;
			3857: outdata = 32'd61679;
			3858: outdata = 32'd61678;
			3859: outdata = 32'd61677;
			3860: outdata = 32'd61676;
			3861: outdata = 32'd61675;
			3862: outdata = 32'd61674;
			3863: outdata = 32'd61673;
			3864: outdata = 32'd61672;
			3865: outdata = 32'd61671;
			3866: outdata = 32'd61670;
			3867: outdata = 32'd61669;
			3868: outdata = 32'd61668;
			3869: outdata = 32'd61667;
			3870: outdata = 32'd61666;
			3871: outdata = 32'd61665;
			3872: outdata = 32'd61664;
			3873: outdata = 32'd61663;
			3874: outdata = 32'd61662;
			3875: outdata = 32'd61661;
			3876: outdata = 32'd61660;
			3877: outdata = 32'd61659;
			3878: outdata = 32'd61658;
			3879: outdata = 32'd61657;
			3880: outdata = 32'd61656;
			3881: outdata = 32'd61655;
			3882: outdata = 32'd61654;
			3883: outdata = 32'd61653;
			3884: outdata = 32'd61652;
			3885: outdata = 32'd61651;
			3886: outdata = 32'd61650;
			3887: outdata = 32'd61649;
			3888: outdata = 32'd61648;
			3889: outdata = 32'd61647;
			3890: outdata = 32'd61646;
			3891: outdata = 32'd61645;
			3892: outdata = 32'd61644;
			3893: outdata = 32'd61643;
			3894: outdata = 32'd61642;
			3895: outdata = 32'd61641;
			3896: outdata = 32'd61640;
			3897: outdata = 32'd61639;
			3898: outdata = 32'd61638;
			3899: outdata = 32'd61637;
			3900: outdata = 32'd61636;
			3901: outdata = 32'd61635;
			3902: outdata = 32'd61634;
			3903: outdata = 32'd61633;
			3904: outdata = 32'd61632;
			3905: outdata = 32'd61631;
			3906: outdata = 32'd61630;
			3907: outdata = 32'd61629;
			3908: outdata = 32'd61628;
			3909: outdata = 32'd61627;
			3910: outdata = 32'd61626;
			3911: outdata = 32'd61625;
			3912: outdata = 32'd61624;
			3913: outdata = 32'd61623;
			3914: outdata = 32'd61622;
			3915: outdata = 32'd61621;
			3916: outdata = 32'd61620;
			3917: outdata = 32'd61619;
			3918: outdata = 32'd61618;
			3919: outdata = 32'd61617;
			3920: outdata = 32'd61616;
			3921: outdata = 32'd61615;
			3922: outdata = 32'd61614;
			3923: outdata = 32'd61613;
			3924: outdata = 32'd61612;
			3925: outdata = 32'd61611;
			3926: outdata = 32'd61610;
			3927: outdata = 32'd61609;
			3928: outdata = 32'd61608;
			3929: outdata = 32'd61607;
			3930: outdata = 32'd61606;
			3931: outdata = 32'd61605;
			3932: outdata = 32'd61604;
			3933: outdata = 32'd61603;
			3934: outdata = 32'd61602;
			3935: outdata = 32'd61601;
			3936: outdata = 32'd61600;
			3937: outdata = 32'd61599;
			3938: outdata = 32'd61598;
			3939: outdata = 32'd61597;
			3940: outdata = 32'd61596;
			3941: outdata = 32'd61595;
			3942: outdata = 32'd61594;
			3943: outdata = 32'd61593;
			3944: outdata = 32'd61592;
			3945: outdata = 32'd61591;
			3946: outdata = 32'd61590;
			3947: outdata = 32'd61589;
			3948: outdata = 32'd61588;
			3949: outdata = 32'd61587;
			3950: outdata = 32'd61586;
			3951: outdata = 32'd61585;
			3952: outdata = 32'd61584;
			3953: outdata = 32'd61583;
			3954: outdata = 32'd61582;
			3955: outdata = 32'd61581;
			3956: outdata = 32'd61580;
			3957: outdata = 32'd61579;
			3958: outdata = 32'd61578;
			3959: outdata = 32'd61577;
			3960: outdata = 32'd61576;
			3961: outdata = 32'd61575;
			3962: outdata = 32'd61574;
			3963: outdata = 32'd61573;
			3964: outdata = 32'd61572;
			3965: outdata = 32'd61571;
			3966: outdata = 32'd61570;
			3967: outdata = 32'd61569;
			3968: outdata = 32'd61568;
			3969: outdata = 32'd61567;
			3970: outdata = 32'd61566;
			3971: outdata = 32'd61565;
			3972: outdata = 32'd61564;
			3973: outdata = 32'd61563;
			3974: outdata = 32'd61562;
			3975: outdata = 32'd61561;
			3976: outdata = 32'd61560;
			3977: outdata = 32'd61559;
			3978: outdata = 32'd61558;
			3979: outdata = 32'd61557;
			3980: outdata = 32'd61556;
			3981: outdata = 32'd61555;
			3982: outdata = 32'd61554;
			3983: outdata = 32'd61553;
			3984: outdata = 32'd61552;
			3985: outdata = 32'd61551;
			3986: outdata = 32'd61550;
			3987: outdata = 32'd61549;
			3988: outdata = 32'd61548;
			3989: outdata = 32'd61547;
			3990: outdata = 32'd61546;
			3991: outdata = 32'd61545;
			3992: outdata = 32'd61544;
			3993: outdata = 32'd61543;
			3994: outdata = 32'd61542;
			3995: outdata = 32'd61541;
			3996: outdata = 32'd61540;
			3997: outdata = 32'd61539;
			3998: outdata = 32'd61538;
			3999: outdata = 32'd61537;
			4000: outdata = 32'd61536;
			4001: outdata = 32'd61535;
			4002: outdata = 32'd61534;
			4003: outdata = 32'd61533;
			4004: outdata = 32'd61532;
			4005: outdata = 32'd61531;
			4006: outdata = 32'd61530;
			4007: outdata = 32'd61529;
			4008: outdata = 32'd61528;
			4009: outdata = 32'd61527;
			4010: outdata = 32'd61526;
			4011: outdata = 32'd61525;
			4012: outdata = 32'd61524;
			4013: outdata = 32'd61523;
			4014: outdata = 32'd61522;
			4015: outdata = 32'd61521;
			4016: outdata = 32'd61520;
			4017: outdata = 32'd61519;
			4018: outdata = 32'd61518;
			4019: outdata = 32'd61517;
			4020: outdata = 32'd61516;
			4021: outdata = 32'd61515;
			4022: outdata = 32'd61514;
			4023: outdata = 32'd61513;
			4024: outdata = 32'd61512;
			4025: outdata = 32'd61511;
			4026: outdata = 32'd61510;
			4027: outdata = 32'd61509;
			4028: outdata = 32'd61508;
			4029: outdata = 32'd61507;
			4030: outdata = 32'd61506;
			4031: outdata = 32'd61505;
			4032: outdata = 32'd61504;
			4033: outdata = 32'd61503;
			4034: outdata = 32'd61502;
			4035: outdata = 32'd61501;
			4036: outdata = 32'd61500;
			4037: outdata = 32'd61499;
			4038: outdata = 32'd61498;
			4039: outdata = 32'd61497;
			4040: outdata = 32'd61496;
			4041: outdata = 32'd61495;
			4042: outdata = 32'd61494;
			4043: outdata = 32'd61493;
			4044: outdata = 32'd61492;
			4045: outdata = 32'd61491;
			4046: outdata = 32'd61490;
			4047: outdata = 32'd61489;
			4048: outdata = 32'd61488;
			4049: outdata = 32'd61487;
			4050: outdata = 32'd61486;
			4051: outdata = 32'd61485;
			4052: outdata = 32'd61484;
			4053: outdata = 32'd61483;
			4054: outdata = 32'd61482;
			4055: outdata = 32'd61481;
			4056: outdata = 32'd61480;
			4057: outdata = 32'd61479;
			4058: outdata = 32'd61478;
			4059: outdata = 32'd61477;
			4060: outdata = 32'd61476;
			4061: outdata = 32'd61475;
			4062: outdata = 32'd61474;
			4063: outdata = 32'd61473;
			4064: outdata = 32'd61472;
			4065: outdata = 32'd61471;
			4066: outdata = 32'd61470;
			4067: outdata = 32'd61469;
			4068: outdata = 32'd61468;
			4069: outdata = 32'd61467;
			4070: outdata = 32'd61466;
			4071: outdata = 32'd61465;
			4072: outdata = 32'd61464;
			4073: outdata = 32'd61463;
			4074: outdata = 32'd61462;
			4075: outdata = 32'd61461;
			4076: outdata = 32'd61460;
			4077: outdata = 32'd61459;
			4078: outdata = 32'd61458;
			4079: outdata = 32'd61457;
			4080: outdata = 32'd61456;
			4081: outdata = 32'd61455;
			4082: outdata = 32'd61454;
			4083: outdata = 32'd61453;
			4084: outdata = 32'd61452;
			4085: outdata = 32'd61451;
			4086: outdata = 32'd61450;
			4087: outdata = 32'd61449;
			4088: outdata = 32'd61448;
			4089: outdata = 32'd61447;
			4090: outdata = 32'd61446;
			4091: outdata = 32'd61445;
			4092: outdata = 32'd61444;
			4093: outdata = 32'd61443;
			4094: outdata = 32'd61442;
			4095: outdata = 32'd61441;
			4096: outdata = 32'd61440;
			4097: outdata = 32'd61439;
			4098: outdata = 32'd61438;
			4099: outdata = 32'd61437;
			4100: outdata = 32'd61436;
			4101: outdata = 32'd61435;
			4102: outdata = 32'd61434;
			4103: outdata = 32'd61433;
			4104: outdata = 32'd61432;
			4105: outdata = 32'd61431;
			4106: outdata = 32'd61430;
			4107: outdata = 32'd61429;
			4108: outdata = 32'd61428;
			4109: outdata = 32'd61427;
			4110: outdata = 32'd61426;
			4111: outdata = 32'd61425;
			4112: outdata = 32'd61424;
			4113: outdata = 32'd61423;
			4114: outdata = 32'd61422;
			4115: outdata = 32'd61421;
			4116: outdata = 32'd61420;
			4117: outdata = 32'd61419;
			4118: outdata = 32'd61418;
			4119: outdata = 32'd61417;
			4120: outdata = 32'd61416;
			4121: outdata = 32'd61415;
			4122: outdata = 32'd61414;
			4123: outdata = 32'd61413;
			4124: outdata = 32'd61412;
			4125: outdata = 32'd61411;
			4126: outdata = 32'd61410;
			4127: outdata = 32'd61409;
			4128: outdata = 32'd61408;
			4129: outdata = 32'd61407;
			4130: outdata = 32'd61406;
			4131: outdata = 32'd61405;
			4132: outdata = 32'd61404;
			4133: outdata = 32'd61403;
			4134: outdata = 32'd61402;
			4135: outdata = 32'd61401;
			4136: outdata = 32'd61400;
			4137: outdata = 32'd61399;
			4138: outdata = 32'd61398;
			4139: outdata = 32'd61397;
			4140: outdata = 32'd61396;
			4141: outdata = 32'd61395;
			4142: outdata = 32'd61394;
			4143: outdata = 32'd61393;
			4144: outdata = 32'd61392;
			4145: outdata = 32'd61391;
			4146: outdata = 32'd61390;
			4147: outdata = 32'd61389;
			4148: outdata = 32'd61388;
			4149: outdata = 32'd61387;
			4150: outdata = 32'd61386;
			4151: outdata = 32'd61385;
			4152: outdata = 32'd61384;
			4153: outdata = 32'd61383;
			4154: outdata = 32'd61382;
			4155: outdata = 32'd61381;
			4156: outdata = 32'd61380;
			4157: outdata = 32'd61379;
			4158: outdata = 32'd61378;
			4159: outdata = 32'd61377;
			4160: outdata = 32'd61376;
			4161: outdata = 32'd61375;
			4162: outdata = 32'd61374;
			4163: outdata = 32'd61373;
			4164: outdata = 32'd61372;
			4165: outdata = 32'd61371;
			4166: outdata = 32'd61370;
			4167: outdata = 32'd61369;
			4168: outdata = 32'd61368;
			4169: outdata = 32'd61367;
			4170: outdata = 32'd61366;
			4171: outdata = 32'd61365;
			4172: outdata = 32'd61364;
			4173: outdata = 32'd61363;
			4174: outdata = 32'd61362;
			4175: outdata = 32'd61361;
			4176: outdata = 32'd61360;
			4177: outdata = 32'd61359;
			4178: outdata = 32'd61358;
			4179: outdata = 32'd61357;
			4180: outdata = 32'd61356;
			4181: outdata = 32'd61355;
			4182: outdata = 32'd61354;
			4183: outdata = 32'd61353;
			4184: outdata = 32'd61352;
			4185: outdata = 32'd61351;
			4186: outdata = 32'd61350;
			4187: outdata = 32'd61349;
			4188: outdata = 32'd61348;
			4189: outdata = 32'd61347;
			4190: outdata = 32'd61346;
			4191: outdata = 32'd61345;
			4192: outdata = 32'd61344;
			4193: outdata = 32'd61343;
			4194: outdata = 32'd61342;
			4195: outdata = 32'd61341;
			4196: outdata = 32'd61340;
			4197: outdata = 32'd61339;
			4198: outdata = 32'd61338;
			4199: outdata = 32'd61337;
			4200: outdata = 32'd61336;
			4201: outdata = 32'd61335;
			4202: outdata = 32'd61334;
			4203: outdata = 32'd61333;
			4204: outdata = 32'd61332;
			4205: outdata = 32'd61331;
			4206: outdata = 32'd61330;
			4207: outdata = 32'd61329;
			4208: outdata = 32'd61328;
			4209: outdata = 32'd61327;
			4210: outdata = 32'd61326;
			4211: outdata = 32'd61325;
			4212: outdata = 32'd61324;
			4213: outdata = 32'd61323;
			4214: outdata = 32'd61322;
			4215: outdata = 32'd61321;
			4216: outdata = 32'd61320;
			4217: outdata = 32'd61319;
			4218: outdata = 32'd61318;
			4219: outdata = 32'd61317;
			4220: outdata = 32'd61316;
			4221: outdata = 32'd61315;
			4222: outdata = 32'd61314;
			4223: outdata = 32'd61313;
			4224: outdata = 32'd61312;
			4225: outdata = 32'd61311;
			4226: outdata = 32'd61310;
			4227: outdata = 32'd61309;
			4228: outdata = 32'd61308;
			4229: outdata = 32'd61307;
			4230: outdata = 32'd61306;
			4231: outdata = 32'd61305;
			4232: outdata = 32'd61304;
			4233: outdata = 32'd61303;
			4234: outdata = 32'd61302;
			4235: outdata = 32'd61301;
			4236: outdata = 32'd61300;
			4237: outdata = 32'd61299;
			4238: outdata = 32'd61298;
			4239: outdata = 32'd61297;
			4240: outdata = 32'd61296;
			4241: outdata = 32'd61295;
			4242: outdata = 32'd61294;
			4243: outdata = 32'd61293;
			4244: outdata = 32'd61292;
			4245: outdata = 32'd61291;
			4246: outdata = 32'd61290;
			4247: outdata = 32'd61289;
			4248: outdata = 32'd61288;
			4249: outdata = 32'd61287;
			4250: outdata = 32'd61286;
			4251: outdata = 32'd61285;
			4252: outdata = 32'd61284;
			4253: outdata = 32'd61283;
			4254: outdata = 32'd61282;
			4255: outdata = 32'd61281;
			4256: outdata = 32'd61280;
			4257: outdata = 32'd61279;
			4258: outdata = 32'd61278;
			4259: outdata = 32'd61277;
			4260: outdata = 32'd61276;
			4261: outdata = 32'd61275;
			4262: outdata = 32'd61274;
			4263: outdata = 32'd61273;
			4264: outdata = 32'd61272;
			4265: outdata = 32'd61271;
			4266: outdata = 32'd61270;
			4267: outdata = 32'd61269;
			4268: outdata = 32'd61268;
			4269: outdata = 32'd61267;
			4270: outdata = 32'd61266;
			4271: outdata = 32'd61265;
			4272: outdata = 32'd61264;
			4273: outdata = 32'd61263;
			4274: outdata = 32'd61262;
			4275: outdata = 32'd61261;
			4276: outdata = 32'd61260;
			4277: outdata = 32'd61259;
			4278: outdata = 32'd61258;
			4279: outdata = 32'd61257;
			4280: outdata = 32'd61256;
			4281: outdata = 32'd61255;
			4282: outdata = 32'd61254;
			4283: outdata = 32'd61253;
			4284: outdata = 32'd61252;
			4285: outdata = 32'd61251;
			4286: outdata = 32'd61250;
			4287: outdata = 32'd61249;
			4288: outdata = 32'd61248;
			4289: outdata = 32'd61247;
			4290: outdata = 32'd61246;
			4291: outdata = 32'd61245;
			4292: outdata = 32'd61244;
			4293: outdata = 32'd61243;
			4294: outdata = 32'd61242;
			4295: outdata = 32'd61241;
			4296: outdata = 32'd61240;
			4297: outdata = 32'd61239;
			4298: outdata = 32'd61238;
			4299: outdata = 32'd61237;
			4300: outdata = 32'd61236;
			4301: outdata = 32'd61235;
			4302: outdata = 32'd61234;
			4303: outdata = 32'd61233;
			4304: outdata = 32'd61232;
			4305: outdata = 32'd61231;
			4306: outdata = 32'd61230;
			4307: outdata = 32'd61229;
			4308: outdata = 32'd61228;
			4309: outdata = 32'd61227;
			4310: outdata = 32'd61226;
			4311: outdata = 32'd61225;
			4312: outdata = 32'd61224;
			4313: outdata = 32'd61223;
			4314: outdata = 32'd61222;
			4315: outdata = 32'd61221;
			4316: outdata = 32'd61220;
			4317: outdata = 32'd61219;
			4318: outdata = 32'd61218;
			4319: outdata = 32'd61217;
			4320: outdata = 32'd61216;
			4321: outdata = 32'd61215;
			4322: outdata = 32'd61214;
			4323: outdata = 32'd61213;
			4324: outdata = 32'd61212;
			4325: outdata = 32'd61211;
			4326: outdata = 32'd61210;
			4327: outdata = 32'd61209;
			4328: outdata = 32'd61208;
			4329: outdata = 32'd61207;
			4330: outdata = 32'd61206;
			4331: outdata = 32'd61205;
			4332: outdata = 32'd61204;
			4333: outdata = 32'd61203;
			4334: outdata = 32'd61202;
			4335: outdata = 32'd61201;
			4336: outdata = 32'd61200;
			4337: outdata = 32'd61199;
			4338: outdata = 32'd61198;
			4339: outdata = 32'd61197;
			4340: outdata = 32'd61196;
			4341: outdata = 32'd61195;
			4342: outdata = 32'd61194;
			4343: outdata = 32'd61193;
			4344: outdata = 32'd61192;
			4345: outdata = 32'd61191;
			4346: outdata = 32'd61190;
			4347: outdata = 32'd61189;
			4348: outdata = 32'd61188;
			4349: outdata = 32'd61187;
			4350: outdata = 32'd61186;
			4351: outdata = 32'd61185;
			4352: outdata = 32'd61184;
			4353: outdata = 32'd61183;
			4354: outdata = 32'd61182;
			4355: outdata = 32'd61181;
			4356: outdata = 32'd61180;
			4357: outdata = 32'd61179;
			4358: outdata = 32'd61178;
			4359: outdata = 32'd61177;
			4360: outdata = 32'd61176;
			4361: outdata = 32'd61175;
			4362: outdata = 32'd61174;
			4363: outdata = 32'd61173;
			4364: outdata = 32'd61172;
			4365: outdata = 32'd61171;
			4366: outdata = 32'd61170;
			4367: outdata = 32'd61169;
			4368: outdata = 32'd61168;
			4369: outdata = 32'd61167;
			4370: outdata = 32'd61166;
			4371: outdata = 32'd61165;
			4372: outdata = 32'd61164;
			4373: outdata = 32'd61163;
			4374: outdata = 32'd61162;
			4375: outdata = 32'd61161;
			4376: outdata = 32'd61160;
			4377: outdata = 32'd61159;
			4378: outdata = 32'd61158;
			4379: outdata = 32'd61157;
			4380: outdata = 32'd61156;
			4381: outdata = 32'd61155;
			4382: outdata = 32'd61154;
			4383: outdata = 32'd61153;
			4384: outdata = 32'd61152;
			4385: outdata = 32'd61151;
			4386: outdata = 32'd61150;
			4387: outdata = 32'd61149;
			4388: outdata = 32'd61148;
			4389: outdata = 32'd61147;
			4390: outdata = 32'd61146;
			4391: outdata = 32'd61145;
			4392: outdata = 32'd61144;
			4393: outdata = 32'd61143;
			4394: outdata = 32'd61142;
			4395: outdata = 32'd61141;
			4396: outdata = 32'd61140;
			4397: outdata = 32'd61139;
			4398: outdata = 32'd61138;
			4399: outdata = 32'd61137;
			4400: outdata = 32'd61136;
			4401: outdata = 32'd61135;
			4402: outdata = 32'd61134;
			4403: outdata = 32'd61133;
			4404: outdata = 32'd61132;
			4405: outdata = 32'd61131;
			4406: outdata = 32'd61130;
			4407: outdata = 32'd61129;
			4408: outdata = 32'd61128;
			4409: outdata = 32'd61127;
			4410: outdata = 32'd61126;
			4411: outdata = 32'd61125;
			4412: outdata = 32'd61124;
			4413: outdata = 32'd61123;
			4414: outdata = 32'd61122;
			4415: outdata = 32'd61121;
			4416: outdata = 32'd61120;
			4417: outdata = 32'd61119;
			4418: outdata = 32'd61118;
			4419: outdata = 32'd61117;
			4420: outdata = 32'd61116;
			4421: outdata = 32'd61115;
			4422: outdata = 32'd61114;
			4423: outdata = 32'd61113;
			4424: outdata = 32'd61112;
			4425: outdata = 32'd61111;
			4426: outdata = 32'd61110;
			4427: outdata = 32'd61109;
			4428: outdata = 32'd61108;
			4429: outdata = 32'd61107;
			4430: outdata = 32'd61106;
			4431: outdata = 32'd61105;
			4432: outdata = 32'd61104;
			4433: outdata = 32'd61103;
			4434: outdata = 32'd61102;
			4435: outdata = 32'd61101;
			4436: outdata = 32'd61100;
			4437: outdata = 32'd61099;
			4438: outdata = 32'd61098;
			4439: outdata = 32'd61097;
			4440: outdata = 32'd61096;
			4441: outdata = 32'd61095;
			4442: outdata = 32'd61094;
			4443: outdata = 32'd61093;
			4444: outdata = 32'd61092;
			4445: outdata = 32'd61091;
			4446: outdata = 32'd61090;
			4447: outdata = 32'd61089;
			4448: outdata = 32'd61088;
			4449: outdata = 32'd61087;
			4450: outdata = 32'd61086;
			4451: outdata = 32'd61085;
			4452: outdata = 32'd61084;
			4453: outdata = 32'd61083;
			4454: outdata = 32'd61082;
			4455: outdata = 32'd61081;
			4456: outdata = 32'd61080;
			4457: outdata = 32'd61079;
			4458: outdata = 32'd61078;
			4459: outdata = 32'd61077;
			4460: outdata = 32'd61076;
			4461: outdata = 32'd61075;
			4462: outdata = 32'd61074;
			4463: outdata = 32'd61073;
			4464: outdata = 32'd61072;
			4465: outdata = 32'd61071;
			4466: outdata = 32'd61070;
			4467: outdata = 32'd61069;
			4468: outdata = 32'd61068;
			4469: outdata = 32'd61067;
			4470: outdata = 32'd61066;
			4471: outdata = 32'd61065;
			4472: outdata = 32'd61064;
			4473: outdata = 32'd61063;
			4474: outdata = 32'd61062;
			4475: outdata = 32'd61061;
			4476: outdata = 32'd61060;
			4477: outdata = 32'd61059;
			4478: outdata = 32'd61058;
			4479: outdata = 32'd61057;
			4480: outdata = 32'd61056;
			4481: outdata = 32'd61055;
			4482: outdata = 32'd61054;
			4483: outdata = 32'd61053;
			4484: outdata = 32'd61052;
			4485: outdata = 32'd61051;
			4486: outdata = 32'd61050;
			4487: outdata = 32'd61049;
			4488: outdata = 32'd61048;
			4489: outdata = 32'd61047;
			4490: outdata = 32'd61046;
			4491: outdata = 32'd61045;
			4492: outdata = 32'd61044;
			4493: outdata = 32'd61043;
			4494: outdata = 32'd61042;
			4495: outdata = 32'd61041;
			4496: outdata = 32'd61040;
			4497: outdata = 32'd61039;
			4498: outdata = 32'd61038;
			4499: outdata = 32'd61037;
			4500: outdata = 32'd61036;
			4501: outdata = 32'd61035;
			4502: outdata = 32'd61034;
			4503: outdata = 32'd61033;
			4504: outdata = 32'd61032;
			4505: outdata = 32'd61031;
			4506: outdata = 32'd61030;
			4507: outdata = 32'd61029;
			4508: outdata = 32'd61028;
			4509: outdata = 32'd61027;
			4510: outdata = 32'd61026;
			4511: outdata = 32'd61025;
			4512: outdata = 32'd61024;
			4513: outdata = 32'd61023;
			4514: outdata = 32'd61022;
			4515: outdata = 32'd61021;
			4516: outdata = 32'd61020;
			4517: outdata = 32'd61019;
			4518: outdata = 32'd61018;
			4519: outdata = 32'd61017;
			4520: outdata = 32'd61016;
			4521: outdata = 32'd61015;
			4522: outdata = 32'd61014;
			4523: outdata = 32'd61013;
			4524: outdata = 32'd61012;
			4525: outdata = 32'd61011;
			4526: outdata = 32'd61010;
			4527: outdata = 32'd61009;
			4528: outdata = 32'd61008;
			4529: outdata = 32'd61007;
			4530: outdata = 32'd61006;
			4531: outdata = 32'd61005;
			4532: outdata = 32'd61004;
			4533: outdata = 32'd61003;
			4534: outdata = 32'd61002;
			4535: outdata = 32'd61001;
			4536: outdata = 32'd61000;
			4537: outdata = 32'd60999;
			4538: outdata = 32'd60998;
			4539: outdata = 32'd60997;
			4540: outdata = 32'd60996;
			4541: outdata = 32'd60995;
			4542: outdata = 32'd60994;
			4543: outdata = 32'd60993;
			4544: outdata = 32'd60992;
			4545: outdata = 32'd60991;
			4546: outdata = 32'd60990;
			4547: outdata = 32'd60989;
			4548: outdata = 32'd60988;
			4549: outdata = 32'd60987;
			4550: outdata = 32'd60986;
			4551: outdata = 32'd60985;
			4552: outdata = 32'd60984;
			4553: outdata = 32'd60983;
			4554: outdata = 32'd60982;
			4555: outdata = 32'd60981;
			4556: outdata = 32'd60980;
			4557: outdata = 32'd60979;
			4558: outdata = 32'd60978;
			4559: outdata = 32'd60977;
			4560: outdata = 32'd60976;
			4561: outdata = 32'd60975;
			4562: outdata = 32'd60974;
			4563: outdata = 32'd60973;
			4564: outdata = 32'd60972;
			4565: outdata = 32'd60971;
			4566: outdata = 32'd60970;
			4567: outdata = 32'd60969;
			4568: outdata = 32'd60968;
			4569: outdata = 32'd60967;
			4570: outdata = 32'd60966;
			4571: outdata = 32'd60965;
			4572: outdata = 32'd60964;
			4573: outdata = 32'd60963;
			4574: outdata = 32'd60962;
			4575: outdata = 32'd60961;
			4576: outdata = 32'd60960;
			4577: outdata = 32'd60959;
			4578: outdata = 32'd60958;
			4579: outdata = 32'd60957;
			4580: outdata = 32'd60956;
			4581: outdata = 32'd60955;
			4582: outdata = 32'd60954;
			4583: outdata = 32'd60953;
			4584: outdata = 32'd60952;
			4585: outdata = 32'd60951;
			4586: outdata = 32'd60950;
			4587: outdata = 32'd60949;
			4588: outdata = 32'd60948;
			4589: outdata = 32'd60947;
			4590: outdata = 32'd60946;
			4591: outdata = 32'd60945;
			4592: outdata = 32'd60944;
			4593: outdata = 32'd60943;
			4594: outdata = 32'd60942;
			4595: outdata = 32'd60941;
			4596: outdata = 32'd60940;
			4597: outdata = 32'd60939;
			4598: outdata = 32'd60938;
			4599: outdata = 32'd60937;
			4600: outdata = 32'd60936;
			4601: outdata = 32'd60935;
			4602: outdata = 32'd60934;
			4603: outdata = 32'd60933;
			4604: outdata = 32'd60932;
			4605: outdata = 32'd60931;
			4606: outdata = 32'd60930;
			4607: outdata = 32'd60929;
			4608: outdata = 32'd60928;
			4609: outdata = 32'd60927;
			4610: outdata = 32'd60926;
			4611: outdata = 32'd60925;
			4612: outdata = 32'd60924;
			4613: outdata = 32'd60923;
			4614: outdata = 32'd60922;
			4615: outdata = 32'd60921;
			4616: outdata = 32'd60920;
			4617: outdata = 32'd60919;
			4618: outdata = 32'd60918;
			4619: outdata = 32'd60917;
			4620: outdata = 32'd60916;
			4621: outdata = 32'd60915;
			4622: outdata = 32'd60914;
			4623: outdata = 32'd60913;
			4624: outdata = 32'd60912;
			4625: outdata = 32'd60911;
			4626: outdata = 32'd60910;
			4627: outdata = 32'd60909;
			4628: outdata = 32'd60908;
			4629: outdata = 32'd60907;
			4630: outdata = 32'd60906;
			4631: outdata = 32'd60905;
			4632: outdata = 32'd60904;
			4633: outdata = 32'd60903;
			4634: outdata = 32'd60902;
			4635: outdata = 32'd60901;
			4636: outdata = 32'd60900;
			4637: outdata = 32'd60899;
			4638: outdata = 32'd60898;
			4639: outdata = 32'd60897;
			4640: outdata = 32'd60896;
			4641: outdata = 32'd60895;
			4642: outdata = 32'd60894;
			4643: outdata = 32'd60893;
			4644: outdata = 32'd60892;
			4645: outdata = 32'd60891;
			4646: outdata = 32'd60890;
			4647: outdata = 32'd60889;
			4648: outdata = 32'd60888;
			4649: outdata = 32'd60887;
			4650: outdata = 32'd60886;
			4651: outdata = 32'd60885;
			4652: outdata = 32'd60884;
			4653: outdata = 32'd60883;
			4654: outdata = 32'd60882;
			4655: outdata = 32'd60881;
			4656: outdata = 32'd60880;
			4657: outdata = 32'd60879;
			4658: outdata = 32'd60878;
			4659: outdata = 32'd60877;
			4660: outdata = 32'd60876;
			4661: outdata = 32'd60875;
			4662: outdata = 32'd60874;
			4663: outdata = 32'd60873;
			4664: outdata = 32'd60872;
			4665: outdata = 32'd60871;
			4666: outdata = 32'd60870;
			4667: outdata = 32'd60869;
			4668: outdata = 32'd60868;
			4669: outdata = 32'd60867;
			4670: outdata = 32'd60866;
			4671: outdata = 32'd60865;
			4672: outdata = 32'd60864;
			4673: outdata = 32'd60863;
			4674: outdata = 32'd60862;
			4675: outdata = 32'd60861;
			4676: outdata = 32'd60860;
			4677: outdata = 32'd60859;
			4678: outdata = 32'd60858;
			4679: outdata = 32'd60857;
			4680: outdata = 32'd60856;
			4681: outdata = 32'd60855;
			4682: outdata = 32'd60854;
			4683: outdata = 32'd60853;
			4684: outdata = 32'd60852;
			4685: outdata = 32'd60851;
			4686: outdata = 32'd60850;
			4687: outdata = 32'd60849;
			4688: outdata = 32'd60848;
			4689: outdata = 32'd60847;
			4690: outdata = 32'd60846;
			4691: outdata = 32'd60845;
			4692: outdata = 32'd60844;
			4693: outdata = 32'd60843;
			4694: outdata = 32'd60842;
			4695: outdata = 32'd60841;
			4696: outdata = 32'd60840;
			4697: outdata = 32'd60839;
			4698: outdata = 32'd60838;
			4699: outdata = 32'd60837;
			4700: outdata = 32'd60836;
			4701: outdata = 32'd60835;
			4702: outdata = 32'd60834;
			4703: outdata = 32'd60833;
			4704: outdata = 32'd60832;
			4705: outdata = 32'd60831;
			4706: outdata = 32'd60830;
			4707: outdata = 32'd60829;
			4708: outdata = 32'd60828;
			4709: outdata = 32'd60827;
			4710: outdata = 32'd60826;
			4711: outdata = 32'd60825;
			4712: outdata = 32'd60824;
			4713: outdata = 32'd60823;
			4714: outdata = 32'd60822;
			4715: outdata = 32'd60821;
			4716: outdata = 32'd60820;
			4717: outdata = 32'd60819;
			4718: outdata = 32'd60818;
			4719: outdata = 32'd60817;
			4720: outdata = 32'd60816;
			4721: outdata = 32'd60815;
			4722: outdata = 32'd60814;
			4723: outdata = 32'd60813;
			4724: outdata = 32'd60812;
			4725: outdata = 32'd60811;
			4726: outdata = 32'd60810;
			4727: outdata = 32'd60809;
			4728: outdata = 32'd60808;
			4729: outdata = 32'd60807;
			4730: outdata = 32'd60806;
			4731: outdata = 32'd60805;
			4732: outdata = 32'd60804;
			4733: outdata = 32'd60803;
			4734: outdata = 32'd60802;
			4735: outdata = 32'd60801;
			4736: outdata = 32'd60800;
			4737: outdata = 32'd60799;
			4738: outdata = 32'd60798;
			4739: outdata = 32'd60797;
			4740: outdata = 32'd60796;
			4741: outdata = 32'd60795;
			4742: outdata = 32'd60794;
			4743: outdata = 32'd60793;
			4744: outdata = 32'd60792;
			4745: outdata = 32'd60791;
			4746: outdata = 32'd60790;
			4747: outdata = 32'd60789;
			4748: outdata = 32'd60788;
			4749: outdata = 32'd60787;
			4750: outdata = 32'd60786;
			4751: outdata = 32'd60785;
			4752: outdata = 32'd60784;
			4753: outdata = 32'd60783;
			4754: outdata = 32'd60782;
			4755: outdata = 32'd60781;
			4756: outdata = 32'd60780;
			4757: outdata = 32'd60779;
			4758: outdata = 32'd60778;
			4759: outdata = 32'd60777;
			4760: outdata = 32'd60776;
			4761: outdata = 32'd60775;
			4762: outdata = 32'd60774;
			4763: outdata = 32'd60773;
			4764: outdata = 32'd60772;
			4765: outdata = 32'd60771;
			4766: outdata = 32'd60770;
			4767: outdata = 32'd60769;
			4768: outdata = 32'd60768;
			4769: outdata = 32'd60767;
			4770: outdata = 32'd60766;
			4771: outdata = 32'd60765;
			4772: outdata = 32'd60764;
			4773: outdata = 32'd60763;
			4774: outdata = 32'd60762;
			4775: outdata = 32'd60761;
			4776: outdata = 32'd60760;
			4777: outdata = 32'd60759;
			4778: outdata = 32'd60758;
			4779: outdata = 32'd60757;
			4780: outdata = 32'd60756;
			4781: outdata = 32'd60755;
			4782: outdata = 32'd60754;
			4783: outdata = 32'd60753;
			4784: outdata = 32'd60752;
			4785: outdata = 32'd60751;
			4786: outdata = 32'd60750;
			4787: outdata = 32'd60749;
			4788: outdata = 32'd60748;
			4789: outdata = 32'd60747;
			4790: outdata = 32'd60746;
			4791: outdata = 32'd60745;
			4792: outdata = 32'd60744;
			4793: outdata = 32'd60743;
			4794: outdata = 32'd60742;
			4795: outdata = 32'd60741;
			4796: outdata = 32'd60740;
			4797: outdata = 32'd60739;
			4798: outdata = 32'd60738;
			4799: outdata = 32'd60737;
			4800: outdata = 32'd60736;
			4801: outdata = 32'd60735;
			4802: outdata = 32'd60734;
			4803: outdata = 32'd60733;
			4804: outdata = 32'd60732;
			4805: outdata = 32'd60731;
			4806: outdata = 32'd60730;
			4807: outdata = 32'd60729;
			4808: outdata = 32'd60728;
			4809: outdata = 32'd60727;
			4810: outdata = 32'd60726;
			4811: outdata = 32'd60725;
			4812: outdata = 32'd60724;
			4813: outdata = 32'd60723;
			4814: outdata = 32'd60722;
			4815: outdata = 32'd60721;
			4816: outdata = 32'd60720;
			4817: outdata = 32'd60719;
			4818: outdata = 32'd60718;
			4819: outdata = 32'd60717;
			4820: outdata = 32'd60716;
			4821: outdata = 32'd60715;
			4822: outdata = 32'd60714;
			4823: outdata = 32'd60713;
			4824: outdata = 32'd60712;
			4825: outdata = 32'd60711;
			4826: outdata = 32'd60710;
			4827: outdata = 32'd60709;
			4828: outdata = 32'd60708;
			4829: outdata = 32'd60707;
			4830: outdata = 32'd60706;
			4831: outdata = 32'd60705;
			4832: outdata = 32'd60704;
			4833: outdata = 32'd60703;
			4834: outdata = 32'd60702;
			4835: outdata = 32'd60701;
			4836: outdata = 32'd60700;
			4837: outdata = 32'd60699;
			4838: outdata = 32'd60698;
			4839: outdata = 32'd60697;
			4840: outdata = 32'd60696;
			4841: outdata = 32'd60695;
			4842: outdata = 32'd60694;
			4843: outdata = 32'd60693;
			4844: outdata = 32'd60692;
			4845: outdata = 32'd60691;
			4846: outdata = 32'd60690;
			4847: outdata = 32'd60689;
			4848: outdata = 32'd60688;
			4849: outdata = 32'd60687;
			4850: outdata = 32'd60686;
			4851: outdata = 32'd60685;
			4852: outdata = 32'd60684;
			4853: outdata = 32'd60683;
			4854: outdata = 32'd60682;
			4855: outdata = 32'd60681;
			4856: outdata = 32'd60680;
			4857: outdata = 32'd60679;
			4858: outdata = 32'd60678;
			4859: outdata = 32'd60677;
			4860: outdata = 32'd60676;
			4861: outdata = 32'd60675;
			4862: outdata = 32'd60674;
			4863: outdata = 32'd60673;
			4864: outdata = 32'd60672;
			4865: outdata = 32'd60671;
			4866: outdata = 32'd60670;
			4867: outdata = 32'd60669;
			4868: outdata = 32'd60668;
			4869: outdata = 32'd60667;
			4870: outdata = 32'd60666;
			4871: outdata = 32'd60665;
			4872: outdata = 32'd60664;
			4873: outdata = 32'd60663;
			4874: outdata = 32'd60662;
			4875: outdata = 32'd60661;
			4876: outdata = 32'd60660;
			4877: outdata = 32'd60659;
			4878: outdata = 32'd60658;
			4879: outdata = 32'd60657;
			4880: outdata = 32'd60656;
			4881: outdata = 32'd60655;
			4882: outdata = 32'd60654;
			4883: outdata = 32'd60653;
			4884: outdata = 32'd60652;
			4885: outdata = 32'd60651;
			4886: outdata = 32'd60650;
			4887: outdata = 32'd60649;
			4888: outdata = 32'd60648;
			4889: outdata = 32'd60647;
			4890: outdata = 32'd60646;
			4891: outdata = 32'd60645;
			4892: outdata = 32'd60644;
			4893: outdata = 32'd60643;
			4894: outdata = 32'd60642;
			4895: outdata = 32'd60641;
			4896: outdata = 32'd60640;
			4897: outdata = 32'd60639;
			4898: outdata = 32'd60638;
			4899: outdata = 32'd60637;
			4900: outdata = 32'd60636;
			4901: outdata = 32'd60635;
			4902: outdata = 32'd60634;
			4903: outdata = 32'd60633;
			4904: outdata = 32'd60632;
			4905: outdata = 32'd60631;
			4906: outdata = 32'd60630;
			4907: outdata = 32'd60629;
			4908: outdata = 32'd60628;
			4909: outdata = 32'd60627;
			4910: outdata = 32'd60626;
			4911: outdata = 32'd60625;
			4912: outdata = 32'd60624;
			4913: outdata = 32'd60623;
			4914: outdata = 32'd60622;
			4915: outdata = 32'd60621;
			4916: outdata = 32'd60620;
			4917: outdata = 32'd60619;
			4918: outdata = 32'd60618;
			4919: outdata = 32'd60617;
			4920: outdata = 32'd60616;
			4921: outdata = 32'd60615;
			4922: outdata = 32'd60614;
			4923: outdata = 32'd60613;
			4924: outdata = 32'd60612;
			4925: outdata = 32'd60611;
			4926: outdata = 32'd60610;
			4927: outdata = 32'd60609;
			4928: outdata = 32'd60608;
			4929: outdata = 32'd60607;
			4930: outdata = 32'd60606;
			4931: outdata = 32'd60605;
			4932: outdata = 32'd60604;
			4933: outdata = 32'd60603;
			4934: outdata = 32'd60602;
			4935: outdata = 32'd60601;
			4936: outdata = 32'd60600;
			4937: outdata = 32'd60599;
			4938: outdata = 32'd60598;
			4939: outdata = 32'd60597;
			4940: outdata = 32'd60596;
			4941: outdata = 32'd60595;
			4942: outdata = 32'd60594;
			4943: outdata = 32'd60593;
			4944: outdata = 32'd60592;
			4945: outdata = 32'd60591;
			4946: outdata = 32'd60590;
			4947: outdata = 32'd60589;
			4948: outdata = 32'd60588;
			4949: outdata = 32'd60587;
			4950: outdata = 32'd60586;
			4951: outdata = 32'd60585;
			4952: outdata = 32'd60584;
			4953: outdata = 32'd60583;
			4954: outdata = 32'd60582;
			4955: outdata = 32'd60581;
			4956: outdata = 32'd60580;
			4957: outdata = 32'd60579;
			4958: outdata = 32'd60578;
			4959: outdata = 32'd60577;
			4960: outdata = 32'd60576;
			4961: outdata = 32'd60575;
			4962: outdata = 32'd60574;
			4963: outdata = 32'd60573;
			4964: outdata = 32'd60572;
			4965: outdata = 32'd60571;
			4966: outdata = 32'd60570;
			4967: outdata = 32'd60569;
			4968: outdata = 32'd60568;
			4969: outdata = 32'd60567;
			4970: outdata = 32'd60566;
			4971: outdata = 32'd60565;
			4972: outdata = 32'd60564;
			4973: outdata = 32'd60563;
			4974: outdata = 32'd60562;
			4975: outdata = 32'd60561;
			4976: outdata = 32'd60560;
			4977: outdata = 32'd60559;
			4978: outdata = 32'd60558;
			4979: outdata = 32'd60557;
			4980: outdata = 32'd60556;
			4981: outdata = 32'd60555;
			4982: outdata = 32'd60554;
			4983: outdata = 32'd60553;
			4984: outdata = 32'd60552;
			4985: outdata = 32'd60551;
			4986: outdata = 32'd60550;
			4987: outdata = 32'd60549;
			4988: outdata = 32'd60548;
			4989: outdata = 32'd60547;
			4990: outdata = 32'd60546;
			4991: outdata = 32'd60545;
			4992: outdata = 32'd60544;
			4993: outdata = 32'd60543;
			4994: outdata = 32'd60542;
			4995: outdata = 32'd60541;
			4996: outdata = 32'd60540;
			4997: outdata = 32'd60539;
			4998: outdata = 32'd60538;
			4999: outdata = 32'd60537;
			5000: outdata = 32'd60536;
			5001: outdata = 32'd60535;
			5002: outdata = 32'd60534;
			5003: outdata = 32'd60533;
			5004: outdata = 32'd60532;
			5005: outdata = 32'd60531;
			5006: outdata = 32'd60530;
			5007: outdata = 32'd60529;
			5008: outdata = 32'd60528;
			5009: outdata = 32'd60527;
			5010: outdata = 32'd60526;
			5011: outdata = 32'd60525;
			5012: outdata = 32'd60524;
			5013: outdata = 32'd60523;
			5014: outdata = 32'd60522;
			5015: outdata = 32'd60521;
			5016: outdata = 32'd60520;
			5017: outdata = 32'd60519;
			5018: outdata = 32'd60518;
			5019: outdata = 32'd60517;
			5020: outdata = 32'd60516;
			5021: outdata = 32'd60515;
			5022: outdata = 32'd60514;
			5023: outdata = 32'd60513;
			5024: outdata = 32'd60512;
			5025: outdata = 32'd60511;
			5026: outdata = 32'd60510;
			5027: outdata = 32'd60509;
			5028: outdata = 32'd60508;
			5029: outdata = 32'd60507;
			5030: outdata = 32'd60506;
			5031: outdata = 32'd60505;
			5032: outdata = 32'd60504;
			5033: outdata = 32'd60503;
			5034: outdata = 32'd60502;
			5035: outdata = 32'd60501;
			5036: outdata = 32'd60500;
			5037: outdata = 32'd60499;
			5038: outdata = 32'd60498;
			5039: outdata = 32'd60497;
			5040: outdata = 32'd60496;
			5041: outdata = 32'd60495;
			5042: outdata = 32'd60494;
			5043: outdata = 32'd60493;
			5044: outdata = 32'd60492;
			5045: outdata = 32'd60491;
			5046: outdata = 32'd60490;
			5047: outdata = 32'd60489;
			5048: outdata = 32'd60488;
			5049: outdata = 32'd60487;
			5050: outdata = 32'd60486;
			5051: outdata = 32'd60485;
			5052: outdata = 32'd60484;
			5053: outdata = 32'd60483;
			5054: outdata = 32'd60482;
			5055: outdata = 32'd60481;
			5056: outdata = 32'd60480;
			5057: outdata = 32'd60479;
			5058: outdata = 32'd60478;
			5059: outdata = 32'd60477;
			5060: outdata = 32'd60476;
			5061: outdata = 32'd60475;
			5062: outdata = 32'd60474;
			5063: outdata = 32'd60473;
			5064: outdata = 32'd60472;
			5065: outdata = 32'd60471;
			5066: outdata = 32'd60470;
			5067: outdata = 32'd60469;
			5068: outdata = 32'd60468;
			5069: outdata = 32'd60467;
			5070: outdata = 32'd60466;
			5071: outdata = 32'd60465;
			5072: outdata = 32'd60464;
			5073: outdata = 32'd60463;
			5074: outdata = 32'd60462;
			5075: outdata = 32'd60461;
			5076: outdata = 32'd60460;
			5077: outdata = 32'd60459;
			5078: outdata = 32'd60458;
			5079: outdata = 32'd60457;
			5080: outdata = 32'd60456;
			5081: outdata = 32'd60455;
			5082: outdata = 32'd60454;
			5083: outdata = 32'd60453;
			5084: outdata = 32'd60452;
			5085: outdata = 32'd60451;
			5086: outdata = 32'd60450;
			5087: outdata = 32'd60449;
			5088: outdata = 32'd60448;
			5089: outdata = 32'd60447;
			5090: outdata = 32'd60446;
			5091: outdata = 32'd60445;
			5092: outdata = 32'd60444;
			5093: outdata = 32'd60443;
			5094: outdata = 32'd60442;
			5095: outdata = 32'd60441;
			5096: outdata = 32'd60440;
			5097: outdata = 32'd60439;
			5098: outdata = 32'd60438;
			5099: outdata = 32'd60437;
			5100: outdata = 32'd60436;
			5101: outdata = 32'd60435;
			5102: outdata = 32'd60434;
			5103: outdata = 32'd60433;
			5104: outdata = 32'd60432;
			5105: outdata = 32'd60431;
			5106: outdata = 32'd60430;
			5107: outdata = 32'd60429;
			5108: outdata = 32'd60428;
			5109: outdata = 32'd60427;
			5110: outdata = 32'd60426;
			5111: outdata = 32'd60425;
			5112: outdata = 32'd60424;
			5113: outdata = 32'd60423;
			5114: outdata = 32'd60422;
			5115: outdata = 32'd60421;
			5116: outdata = 32'd60420;
			5117: outdata = 32'd60419;
			5118: outdata = 32'd60418;
			5119: outdata = 32'd60417;
			5120: outdata = 32'd60416;
			5121: outdata = 32'd60415;
			5122: outdata = 32'd60414;
			5123: outdata = 32'd60413;
			5124: outdata = 32'd60412;
			5125: outdata = 32'd60411;
			5126: outdata = 32'd60410;
			5127: outdata = 32'd60409;
			5128: outdata = 32'd60408;
			5129: outdata = 32'd60407;
			5130: outdata = 32'd60406;
			5131: outdata = 32'd60405;
			5132: outdata = 32'd60404;
			5133: outdata = 32'd60403;
			5134: outdata = 32'd60402;
			5135: outdata = 32'd60401;
			5136: outdata = 32'd60400;
			5137: outdata = 32'd60399;
			5138: outdata = 32'd60398;
			5139: outdata = 32'd60397;
			5140: outdata = 32'd60396;
			5141: outdata = 32'd60395;
			5142: outdata = 32'd60394;
			5143: outdata = 32'd60393;
			5144: outdata = 32'd60392;
			5145: outdata = 32'd60391;
			5146: outdata = 32'd60390;
			5147: outdata = 32'd60389;
			5148: outdata = 32'd60388;
			5149: outdata = 32'd60387;
			5150: outdata = 32'd60386;
			5151: outdata = 32'd60385;
			5152: outdata = 32'd60384;
			5153: outdata = 32'd60383;
			5154: outdata = 32'd60382;
			5155: outdata = 32'd60381;
			5156: outdata = 32'd60380;
			5157: outdata = 32'd60379;
			5158: outdata = 32'd60378;
			5159: outdata = 32'd60377;
			5160: outdata = 32'd60376;
			5161: outdata = 32'd60375;
			5162: outdata = 32'd60374;
			5163: outdata = 32'd60373;
			5164: outdata = 32'd60372;
			5165: outdata = 32'd60371;
			5166: outdata = 32'd60370;
			5167: outdata = 32'd60369;
			5168: outdata = 32'd60368;
			5169: outdata = 32'd60367;
			5170: outdata = 32'd60366;
			5171: outdata = 32'd60365;
			5172: outdata = 32'd60364;
			5173: outdata = 32'd60363;
			5174: outdata = 32'd60362;
			5175: outdata = 32'd60361;
			5176: outdata = 32'd60360;
			5177: outdata = 32'd60359;
			5178: outdata = 32'd60358;
			5179: outdata = 32'd60357;
			5180: outdata = 32'd60356;
			5181: outdata = 32'd60355;
			5182: outdata = 32'd60354;
			5183: outdata = 32'd60353;
			5184: outdata = 32'd60352;
			5185: outdata = 32'd60351;
			5186: outdata = 32'd60350;
			5187: outdata = 32'd60349;
			5188: outdata = 32'd60348;
			5189: outdata = 32'd60347;
			5190: outdata = 32'd60346;
			5191: outdata = 32'd60345;
			5192: outdata = 32'd60344;
			5193: outdata = 32'd60343;
			5194: outdata = 32'd60342;
			5195: outdata = 32'd60341;
			5196: outdata = 32'd60340;
			5197: outdata = 32'd60339;
			5198: outdata = 32'd60338;
			5199: outdata = 32'd60337;
			5200: outdata = 32'd60336;
			5201: outdata = 32'd60335;
			5202: outdata = 32'd60334;
			5203: outdata = 32'd60333;
			5204: outdata = 32'd60332;
			5205: outdata = 32'd60331;
			5206: outdata = 32'd60330;
			5207: outdata = 32'd60329;
			5208: outdata = 32'd60328;
			5209: outdata = 32'd60327;
			5210: outdata = 32'd60326;
			5211: outdata = 32'd60325;
			5212: outdata = 32'd60324;
			5213: outdata = 32'd60323;
			5214: outdata = 32'd60322;
			5215: outdata = 32'd60321;
			5216: outdata = 32'd60320;
			5217: outdata = 32'd60319;
			5218: outdata = 32'd60318;
			5219: outdata = 32'd60317;
			5220: outdata = 32'd60316;
			5221: outdata = 32'd60315;
			5222: outdata = 32'd60314;
			5223: outdata = 32'd60313;
			5224: outdata = 32'd60312;
			5225: outdata = 32'd60311;
			5226: outdata = 32'd60310;
			5227: outdata = 32'd60309;
			5228: outdata = 32'd60308;
			5229: outdata = 32'd60307;
			5230: outdata = 32'd60306;
			5231: outdata = 32'd60305;
			5232: outdata = 32'd60304;
			5233: outdata = 32'd60303;
			5234: outdata = 32'd60302;
			5235: outdata = 32'd60301;
			5236: outdata = 32'd60300;
			5237: outdata = 32'd60299;
			5238: outdata = 32'd60298;
			5239: outdata = 32'd60297;
			5240: outdata = 32'd60296;
			5241: outdata = 32'd60295;
			5242: outdata = 32'd60294;
			5243: outdata = 32'd60293;
			5244: outdata = 32'd60292;
			5245: outdata = 32'd60291;
			5246: outdata = 32'd60290;
			5247: outdata = 32'd60289;
			5248: outdata = 32'd60288;
			5249: outdata = 32'd60287;
			5250: outdata = 32'd60286;
			5251: outdata = 32'd60285;
			5252: outdata = 32'd60284;
			5253: outdata = 32'd60283;
			5254: outdata = 32'd60282;
			5255: outdata = 32'd60281;
			5256: outdata = 32'd60280;
			5257: outdata = 32'd60279;
			5258: outdata = 32'd60278;
			5259: outdata = 32'd60277;
			5260: outdata = 32'd60276;
			5261: outdata = 32'd60275;
			5262: outdata = 32'd60274;
			5263: outdata = 32'd60273;
			5264: outdata = 32'd60272;
			5265: outdata = 32'd60271;
			5266: outdata = 32'd60270;
			5267: outdata = 32'd60269;
			5268: outdata = 32'd60268;
			5269: outdata = 32'd60267;
			5270: outdata = 32'd60266;
			5271: outdata = 32'd60265;
			5272: outdata = 32'd60264;
			5273: outdata = 32'd60263;
			5274: outdata = 32'd60262;
			5275: outdata = 32'd60261;
			5276: outdata = 32'd60260;
			5277: outdata = 32'd60259;
			5278: outdata = 32'd60258;
			5279: outdata = 32'd60257;
			5280: outdata = 32'd60256;
			5281: outdata = 32'd60255;
			5282: outdata = 32'd60254;
			5283: outdata = 32'd60253;
			5284: outdata = 32'd60252;
			5285: outdata = 32'd60251;
			5286: outdata = 32'd60250;
			5287: outdata = 32'd60249;
			5288: outdata = 32'd60248;
			5289: outdata = 32'd60247;
			5290: outdata = 32'd60246;
			5291: outdata = 32'd60245;
			5292: outdata = 32'd60244;
			5293: outdata = 32'd60243;
			5294: outdata = 32'd60242;
			5295: outdata = 32'd60241;
			5296: outdata = 32'd60240;
			5297: outdata = 32'd60239;
			5298: outdata = 32'd60238;
			5299: outdata = 32'd60237;
			5300: outdata = 32'd60236;
			5301: outdata = 32'd60235;
			5302: outdata = 32'd60234;
			5303: outdata = 32'd60233;
			5304: outdata = 32'd60232;
			5305: outdata = 32'd60231;
			5306: outdata = 32'd60230;
			5307: outdata = 32'd60229;
			5308: outdata = 32'd60228;
			5309: outdata = 32'd60227;
			5310: outdata = 32'd60226;
			5311: outdata = 32'd60225;
			5312: outdata = 32'd60224;
			5313: outdata = 32'd60223;
			5314: outdata = 32'd60222;
			5315: outdata = 32'd60221;
			5316: outdata = 32'd60220;
			5317: outdata = 32'd60219;
			5318: outdata = 32'd60218;
			5319: outdata = 32'd60217;
			5320: outdata = 32'd60216;
			5321: outdata = 32'd60215;
			5322: outdata = 32'd60214;
			5323: outdata = 32'd60213;
			5324: outdata = 32'd60212;
			5325: outdata = 32'd60211;
			5326: outdata = 32'd60210;
			5327: outdata = 32'd60209;
			5328: outdata = 32'd60208;
			5329: outdata = 32'd60207;
			5330: outdata = 32'd60206;
			5331: outdata = 32'd60205;
			5332: outdata = 32'd60204;
			5333: outdata = 32'd60203;
			5334: outdata = 32'd60202;
			5335: outdata = 32'd60201;
			5336: outdata = 32'd60200;
			5337: outdata = 32'd60199;
			5338: outdata = 32'd60198;
			5339: outdata = 32'd60197;
			5340: outdata = 32'd60196;
			5341: outdata = 32'd60195;
			5342: outdata = 32'd60194;
			5343: outdata = 32'd60193;
			5344: outdata = 32'd60192;
			5345: outdata = 32'd60191;
			5346: outdata = 32'd60190;
			5347: outdata = 32'd60189;
			5348: outdata = 32'd60188;
			5349: outdata = 32'd60187;
			5350: outdata = 32'd60186;
			5351: outdata = 32'd60185;
			5352: outdata = 32'd60184;
			5353: outdata = 32'd60183;
			5354: outdata = 32'd60182;
			5355: outdata = 32'd60181;
			5356: outdata = 32'd60180;
			5357: outdata = 32'd60179;
			5358: outdata = 32'd60178;
			5359: outdata = 32'd60177;
			5360: outdata = 32'd60176;
			5361: outdata = 32'd60175;
			5362: outdata = 32'd60174;
			5363: outdata = 32'd60173;
			5364: outdata = 32'd60172;
			5365: outdata = 32'd60171;
			5366: outdata = 32'd60170;
			5367: outdata = 32'd60169;
			5368: outdata = 32'd60168;
			5369: outdata = 32'd60167;
			5370: outdata = 32'd60166;
			5371: outdata = 32'd60165;
			5372: outdata = 32'd60164;
			5373: outdata = 32'd60163;
			5374: outdata = 32'd60162;
			5375: outdata = 32'd60161;
			5376: outdata = 32'd60160;
			5377: outdata = 32'd60159;
			5378: outdata = 32'd60158;
			5379: outdata = 32'd60157;
			5380: outdata = 32'd60156;
			5381: outdata = 32'd60155;
			5382: outdata = 32'd60154;
			5383: outdata = 32'd60153;
			5384: outdata = 32'd60152;
			5385: outdata = 32'd60151;
			5386: outdata = 32'd60150;
			5387: outdata = 32'd60149;
			5388: outdata = 32'd60148;
			5389: outdata = 32'd60147;
			5390: outdata = 32'd60146;
			5391: outdata = 32'd60145;
			5392: outdata = 32'd60144;
			5393: outdata = 32'd60143;
			5394: outdata = 32'd60142;
			5395: outdata = 32'd60141;
			5396: outdata = 32'd60140;
			5397: outdata = 32'd60139;
			5398: outdata = 32'd60138;
			5399: outdata = 32'd60137;
			5400: outdata = 32'd60136;
			5401: outdata = 32'd60135;
			5402: outdata = 32'd60134;
			5403: outdata = 32'd60133;
			5404: outdata = 32'd60132;
			5405: outdata = 32'd60131;
			5406: outdata = 32'd60130;
			5407: outdata = 32'd60129;
			5408: outdata = 32'd60128;
			5409: outdata = 32'd60127;
			5410: outdata = 32'd60126;
			5411: outdata = 32'd60125;
			5412: outdata = 32'd60124;
			5413: outdata = 32'd60123;
			5414: outdata = 32'd60122;
			5415: outdata = 32'd60121;
			5416: outdata = 32'd60120;
			5417: outdata = 32'd60119;
			5418: outdata = 32'd60118;
			5419: outdata = 32'd60117;
			5420: outdata = 32'd60116;
			5421: outdata = 32'd60115;
			5422: outdata = 32'd60114;
			5423: outdata = 32'd60113;
			5424: outdata = 32'd60112;
			5425: outdata = 32'd60111;
			5426: outdata = 32'd60110;
			5427: outdata = 32'd60109;
			5428: outdata = 32'd60108;
			5429: outdata = 32'd60107;
			5430: outdata = 32'd60106;
			5431: outdata = 32'd60105;
			5432: outdata = 32'd60104;
			5433: outdata = 32'd60103;
			5434: outdata = 32'd60102;
			5435: outdata = 32'd60101;
			5436: outdata = 32'd60100;
			5437: outdata = 32'd60099;
			5438: outdata = 32'd60098;
			5439: outdata = 32'd60097;
			5440: outdata = 32'd60096;
			5441: outdata = 32'd60095;
			5442: outdata = 32'd60094;
			5443: outdata = 32'd60093;
			5444: outdata = 32'd60092;
			5445: outdata = 32'd60091;
			5446: outdata = 32'd60090;
			5447: outdata = 32'd60089;
			5448: outdata = 32'd60088;
			5449: outdata = 32'd60087;
			5450: outdata = 32'd60086;
			5451: outdata = 32'd60085;
			5452: outdata = 32'd60084;
			5453: outdata = 32'd60083;
			5454: outdata = 32'd60082;
			5455: outdata = 32'd60081;
			5456: outdata = 32'd60080;
			5457: outdata = 32'd60079;
			5458: outdata = 32'd60078;
			5459: outdata = 32'd60077;
			5460: outdata = 32'd60076;
			5461: outdata = 32'd60075;
			5462: outdata = 32'd60074;
			5463: outdata = 32'd60073;
			5464: outdata = 32'd60072;
			5465: outdata = 32'd60071;
			5466: outdata = 32'd60070;
			5467: outdata = 32'd60069;
			5468: outdata = 32'd60068;
			5469: outdata = 32'd60067;
			5470: outdata = 32'd60066;
			5471: outdata = 32'd60065;
			5472: outdata = 32'd60064;
			5473: outdata = 32'd60063;
			5474: outdata = 32'd60062;
			5475: outdata = 32'd60061;
			5476: outdata = 32'd60060;
			5477: outdata = 32'd60059;
			5478: outdata = 32'd60058;
			5479: outdata = 32'd60057;
			5480: outdata = 32'd60056;
			5481: outdata = 32'd60055;
			5482: outdata = 32'd60054;
			5483: outdata = 32'd60053;
			5484: outdata = 32'd60052;
			5485: outdata = 32'd60051;
			5486: outdata = 32'd60050;
			5487: outdata = 32'd60049;
			5488: outdata = 32'd60048;
			5489: outdata = 32'd60047;
			5490: outdata = 32'd60046;
			5491: outdata = 32'd60045;
			5492: outdata = 32'd60044;
			5493: outdata = 32'd60043;
			5494: outdata = 32'd60042;
			5495: outdata = 32'd60041;
			5496: outdata = 32'd60040;
			5497: outdata = 32'd60039;
			5498: outdata = 32'd60038;
			5499: outdata = 32'd60037;
			5500: outdata = 32'd60036;
			5501: outdata = 32'd60035;
			5502: outdata = 32'd60034;
			5503: outdata = 32'd60033;
			5504: outdata = 32'd60032;
			5505: outdata = 32'd60031;
			5506: outdata = 32'd60030;
			5507: outdata = 32'd60029;
			5508: outdata = 32'd60028;
			5509: outdata = 32'd60027;
			5510: outdata = 32'd60026;
			5511: outdata = 32'd60025;
			5512: outdata = 32'd60024;
			5513: outdata = 32'd60023;
			5514: outdata = 32'd60022;
			5515: outdata = 32'd60021;
			5516: outdata = 32'd60020;
			5517: outdata = 32'd60019;
			5518: outdata = 32'd60018;
			5519: outdata = 32'd60017;
			5520: outdata = 32'd60016;
			5521: outdata = 32'd60015;
			5522: outdata = 32'd60014;
			5523: outdata = 32'd60013;
			5524: outdata = 32'd60012;
			5525: outdata = 32'd60011;
			5526: outdata = 32'd60010;
			5527: outdata = 32'd60009;
			5528: outdata = 32'd60008;
			5529: outdata = 32'd60007;
			5530: outdata = 32'd60006;
			5531: outdata = 32'd60005;
			5532: outdata = 32'd60004;
			5533: outdata = 32'd60003;
			5534: outdata = 32'd60002;
			5535: outdata = 32'd60001;
			5536: outdata = 32'd60000;
			5537: outdata = 32'd59999;
			5538: outdata = 32'd59998;
			5539: outdata = 32'd59997;
			5540: outdata = 32'd59996;
			5541: outdata = 32'd59995;
			5542: outdata = 32'd59994;
			5543: outdata = 32'd59993;
			5544: outdata = 32'd59992;
			5545: outdata = 32'd59991;
			5546: outdata = 32'd59990;
			5547: outdata = 32'd59989;
			5548: outdata = 32'd59988;
			5549: outdata = 32'd59987;
			5550: outdata = 32'd59986;
			5551: outdata = 32'd59985;
			5552: outdata = 32'd59984;
			5553: outdata = 32'd59983;
			5554: outdata = 32'd59982;
			5555: outdata = 32'd59981;
			5556: outdata = 32'd59980;
			5557: outdata = 32'd59979;
			5558: outdata = 32'd59978;
			5559: outdata = 32'd59977;
			5560: outdata = 32'd59976;
			5561: outdata = 32'd59975;
			5562: outdata = 32'd59974;
			5563: outdata = 32'd59973;
			5564: outdata = 32'd59972;
			5565: outdata = 32'd59971;
			5566: outdata = 32'd59970;
			5567: outdata = 32'd59969;
			5568: outdata = 32'd59968;
			5569: outdata = 32'd59967;
			5570: outdata = 32'd59966;
			5571: outdata = 32'd59965;
			5572: outdata = 32'd59964;
			5573: outdata = 32'd59963;
			5574: outdata = 32'd59962;
			5575: outdata = 32'd59961;
			5576: outdata = 32'd59960;
			5577: outdata = 32'd59959;
			5578: outdata = 32'd59958;
			5579: outdata = 32'd59957;
			5580: outdata = 32'd59956;
			5581: outdata = 32'd59955;
			5582: outdata = 32'd59954;
			5583: outdata = 32'd59953;
			5584: outdata = 32'd59952;
			5585: outdata = 32'd59951;
			5586: outdata = 32'd59950;
			5587: outdata = 32'd59949;
			5588: outdata = 32'd59948;
			5589: outdata = 32'd59947;
			5590: outdata = 32'd59946;
			5591: outdata = 32'd59945;
			5592: outdata = 32'd59944;
			5593: outdata = 32'd59943;
			5594: outdata = 32'd59942;
			5595: outdata = 32'd59941;
			5596: outdata = 32'd59940;
			5597: outdata = 32'd59939;
			5598: outdata = 32'd59938;
			5599: outdata = 32'd59937;
			5600: outdata = 32'd59936;
			5601: outdata = 32'd59935;
			5602: outdata = 32'd59934;
			5603: outdata = 32'd59933;
			5604: outdata = 32'd59932;
			5605: outdata = 32'd59931;
			5606: outdata = 32'd59930;
			5607: outdata = 32'd59929;
			5608: outdata = 32'd59928;
			5609: outdata = 32'd59927;
			5610: outdata = 32'd59926;
			5611: outdata = 32'd59925;
			5612: outdata = 32'd59924;
			5613: outdata = 32'd59923;
			5614: outdata = 32'd59922;
			5615: outdata = 32'd59921;
			5616: outdata = 32'd59920;
			5617: outdata = 32'd59919;
			5618: outdata = 32'd59918;
			5619: outdata = 32'd59917;
			5620: outdata = 32'd59916;
			5621: outdata = 32'd59915;
			5622: outdata = 32'd59914;
			5623: outdata = 32'd59913;
			5624: outdata = 32'd59912;
			5625: outdata = 32'd59911;
			5626: outdata = 32'd59910;
			5627: outdata = 32'd59909;
			5628: outdata = 32'd59908;
			5629: outdata = 32'd59907;
			5630: outdata = 32'd59906;
			5631: outdata = 32'd59905;
			5632: outdata = 32'd59904;
			5633: outdata = 32'd59903;
			5634: outdata = 32'd59902;
			5635: outdata = 32'd59901;
			5636: outdata = 32'd59900;
			5637: outdata = 32'd59899;
			5638: outdata = 32'd59898;
			5639: outdata = 32'd59897;
			5640: outdata = 32'd59896;
			5641: outdata = 32'd59895;
			5642: outdata = 32'd59894;
			5643: outdata = 32'd59893;
			5644: outdata = 32'd59892;
			5645: outdata = 32'd59891;
			5646: outdata = 32'd59890;
			5647: outdata = 32'd59889;
			5648: outdata = 32'd59888;
			5649: outdata = 32'd59887;
			5650: outdata = 32'd59886;
			5651: outdata = 32'd59885;
			5652: outdata = 32'd59884;
			5653: outdata = 32'd59883;
			5654: outdata = 32'd59882;
			5655: outdata = 32'd59881;
			5656: outdata = 32'd59880;
			5657: outdata = 32'd59879;
			5658: outdata = 32'd59878;
			5659: outdata = 32'd59877;
			5660: outdata = 32'd59876;
			5661: outdata = 32'd59875;
			5662: outdata = 32'd59874;
			5663: outdata = 32'd59873;
			5664: outdata = 32'd59872;
			5665: outdata = 32'd59871;
			5666: outdata = 32'd59870;
			5667: outdata = 32'd59869;
			5668: outdata = 32'd59868;
			5669: outdata = 32'd59867;
			5670: outdata = 32'd59866;
			5671: outdata = 32'd59865;
			5672: outdata = 32'd59864;
			5673: outdata = 32'd59863;
			5674: outdata = 32'd59862;
			5675: outdata = 32'd59861;
			5676: outdata = 32'd59860;
			5677: outdata = 32'd59859;
			5678: outdata = 32'd59858;
			5679: outdata = 32'd59857;
			5680: outdata = 32'd59856;
			5681: outdata = 32'd59855;
			5682: outdata = 32'd59854;
			5683: outdata = 32'd59853;
			5684: outdata = 32'd59852;
			5685: outdata = 32'd59851;
			5686: outdata = 32'd59850;
			5687: outdata = 32'd59849;
			5688: outdata = 32'd59848;
			5689: outdata = 32'd59847;
			5690: outdata = 32'd59846;
			5691: outdata = 32'd59845;
			5692: outdata = 32'd59844;
			5693: outdata = 32'd59843;
			5694: outdata = 32'd59842;
			5695: outdata = 32'd59841;
			5696: outdata = 32'd59840;
			5697: outdata = 32'd59839;
			5698: outdata = 32'd59838;
			5699: outdata = 32'd59837;
			5700: outdata = 32'd59836;
			5701: outdata = 32'd59835;
			5702: outdata = 32'd59834;
			5703: outdata = 32'd59833;
			5704: outdata = 32'd59832;
			5705: outdata = 32'd59831;
			5706: outdata = 32'd59830;
			5707: outdata = 32'd59829;
			5708: outdata = 32'd59828;
			5709: outdata = 32'd59827;
			5710: outdata = 32'd59826;
			5711: outdata = 32'd59825;
			5712: outdata = 32'd59824;
			5713: outdata = 32'd59823;
			5714: outdata = 32'd59822;
			5715: outdata = 32'd59821;
			5716: outdata = 32'd59820;
			5717: outdata = 32'd59819;
			5718: outdata = 32'd59818;
			5719: outdata = 32'd59817;
			5720: outdata = 32'd59816;
			5721: outdata = 32'd59815;
			5722: outdata = 32'd59814;
			5723: outdata = 32'd59813;
			5724: outdata = 32'd59812;
			5725: outdata = 32'd59811;
			5726: outdata = 32'd59810;
			5727: outdata = 32'd59809;
			5728: outdata = 32'd59808;
			5729: outdata = 32'd59807;
			5730: outdata = 32'd59806;
			5731: outdata = 32'd59805;
			5732: outdata = 32'd59804;
			5733: outdata = 32'd59803;
			5734: outdata = 32'd59802;
			5735: outdata = 32'd59801;
			5736: outdata = 32'd59800;
			5737: outdata = 32'd59799;
			5738: outdata = 32'd59798;
			5739: outdata = 32'd59797;
			5740: outdata = 32'd59796;
			5741: outdata = 32'd59795;
			5742: outdata = 32'd59794;
			5743: outdata = 32'd59793;
			5744: outdata = 32'd59792;
			5745: outdata = 32'd59791;
			5746: outdata = 32'd59790;
			5747: outdata = 32'd59789;
			5748: outdata = 32'd59788;
			5749: outdata = 32'd59787;
			5750: outdata = 32'd59786;
			5751: outdata = 32'd59785;
			5752: outdata = 32'd59784;
			5753: outdata = 32'd59783;
			5754: outdata = 32'd59782;
			5755: outdata = 32'd59781;
			5756: outdata = 32'd59780;
			5757: outdata = 32'd59779;
			5758: outdata = 32'd59778;
			5759: outdata = 32'd59777;
			5760: outdata = 32'd59776;
			5761: outdata = 32'd59775;
			5762: outdata = 32'd59774;
			5763: outdata = 32'd59773;
			5764: outdata = 32'd59772;
			5765: outdata = 32'd59771;
			5766: outdata = 32'd59770;
			5767: outdata = 32'd59769;
			5768: outdata = 32'd59768;
			5769: outdata = 32'd59767;
			5770: outdata = 32'd59766;
			5771: outdata = 32'd59765;
			5772: outdata = 32'd59764;
			5773: outdata = 32'd59763;
			5774: outdata = 32'd59762;
			5775: outdata = 32'd59761;
			5776: outdata = 32'd59760;
			5777: outdata = 32'd59759;
			5778: outdata = 32'd59758;
			5779: outdata = 32'd59757;
			5780: outdata = 32'd59756;
			5781: outdata = 32'd59755;
			5782: outdata = 32'd59754;
			5783: outdata = 32'd59753;
			5784: outdata = 32'd59752;
			5785: outdata = 32'd59751;
			5786: outdata = 32'd59750;
			5787: outdata = 32'd59749;
			5788: outdata = 32'd59748;
			5789: outdata = 32'd59747;
			5790: outdata = 32'd59746;
			5791: outdata = 32'd59745;
			5792: outdata = 32'd59744;
			5793: outdata = 32'd59743;
			5794: outdata = 32'd59742;
			5795: outdata = 32'd59741;
			5796: outdata = 32'd59740;
			5797: outdata = 32'd59739;
			5798: outdata = 32'd59738;
			5799: outdata = 32'd59737;
			5800: outdata = 32'd59736;
			5801: outdata = 32'd59735;
			5802: outdata = 32'd59734;
			5803: outdata = 32'd59733;
			5804: outdata = 32'd59732;
			5805: outdata = 32'd59731;
			5806: outdata = 32'd59730;
			5807: outdata = 32'd59729;
			5808: outdata = 32'd59728;
			5809: outdata = 32'd59727;
			5810: outdata = 32'd59726;
			5811: outdata = 32'd59725;
			5812: outdata = 32'd59724;
			5813: outdata = 32'd59723;
			5814: outdata = 32'd59722;
			5815: outdata = 32'd59721;
			5816: outdata = 32'd59720;
			5817: outdata = 32'd59719;
			5818: outdata = 32'd59718;
			5819: outdata = 32'd59717;
			5820: outdata = 32'd59716;
			5821: outdata = 32'd59715;
			5822: outdata = 32'd59714;
			5823: outdata = 32'd59713;
			5824: outdata = 32'd59712;
			5825: outdata = 32'd59711;
			5826: outdata = 32'd59710;
			5827: outdata = 32'd59709;
			5828: outdata = 32'd59708;
			5829: outdata = 32'd59707;
			5830: outdata = 32'd59706;
			5831: outdata = 32'd59705;
			5832: outdata = 32'd59704;
			5833: outdata = 32'd59703;
			5834: outdata = 32'd59702;
			5835: outdata = 32'd59701;
			5836: outdata = 32'd59700;
			5837: outdata = 32'd59699;
			5838: outdata = 32'd59698;
			5839: outdata = 32'd59697;
			5840: outdata = 32'd59696;
			5841: outdata = 32'd59695;
			5842: outdata = 32'd59694;
			5843: outdata = 32'd59693;
			5844: outdata = 32'd59692;
			5845: outdata = 32'd59691;
			5846: outdata = 32'd59690;
			5847: outdata = 32'd59689;
			5848: outdata = 32'd59688;
			5849: outdata = 32'd59687;
			5850: outdata = 32'd59686;
			5851: outdata = 32'd59685;
			5852: outdata = 32'd59684;
			5853: outdata = 32'd59683;
			5854: outdata = 32'd59682;
			5855: outdata = 32'd59681;
			5856: outdata = 32'd59680;
			5857: outdata = 32'd59679;
			5858: outdata = 32'd59678;
			5859: outdata = 32'd59677;
			5860: outdata = 32'd59676;
			5861: outdata = 32'd59675;
			5862: outdata = 32'd59674;
			5863: outdata = 32'd59673;
			5864: outdata = 32'd59672;
			5865: outdata = 32'd59671;
			5866: outdata = 32'd59670;
			5867: outdata = 32'd59669;
			5868: outdata = 32'd59668;
			5869: outdata = 32'd59667;
			5870: outdata = 32'd59666;
			5871: outdata = 32'd59665;
			5872: outdata = 32'd59664;
			5873: outdata = 32'd59663;
			5874: outdata = 32'd59662;
			5875: outdata = 32'd59661;
			5876: outdata = 32'd59660;
			5877: outdata = 32'd59659;
			5878: outdata = 32'd59658;
			5879: outdata = 32'd59657;
			5880: outdata = 32'd59656;
			5881: outdata = 32'd59655;
			5882: outdata = 32'd59654;
			5883: outdata = 32'd59653;
			5884: outdata = 32'd59652;
			5885: outdata = 32'd59651;
			5886: outdata = 32'd59650;
			5887: outdata = 32'd59649;
			5888: outdata = 32'd59648;
			5889: outdata = 32'd59647;
			5890: outdata = 32'd59646;
			5891: outdata = 32'd59645;
			5892: outdata = 32'd59644;
			5893: outdata = 32'd59643;
			5894: outdata = 32'd59642;
			5895: outdata = 32'd59641;
			5896: outdata = 32'd59640;
			5897: outdata = 32'd59639;
			5898: outdata = 32'd59638;
			5899: outdata = 32'd59637;
			5900: outdata = 32'd59636;
			5901: outdata = 32'd59635;
			5902: outdata = 32'd59634;
			5903: outdata = 32'd59633;
			5904: outdata = 32'd59632;
			5905: outdata = 32'd59631;
			5906: outdata = 32'd59630;
			5907: outdata = 32'd59629;
			5908: outdata = 32'd59628;
			5909: outdata = 32'd59627;
			5910: outdata = 32'd59626;
			5911: outdata = 32'd59625;
			5912: outdata = 32'd59624;
			5913: outdata = 32'd59623;
			5914: outdata = 32'd59622;
			5915: outdata = 32'd59621;
			5916: outdata = 32'd59620;
			5917: outdata = 32'd59619;
			5918: outdata = 32'd59618;
			5919: outdata = 32'd59617;
			5920: outdata = 32'd59616;
			5921: outdata = 32'd59615;
			5922: outdata = 32'd59614;
			5923: outdata = 32'd59613;
			5924: outdata = 32'd59612;
			5925: outdata = 32'd59611;
			5926: outdata = 32'd59610;
			5927: outdata = 32'd59609;
			5928: outdata = 32'd59608;
			5929: outdata = 32'd59607;
			5930: outdata = 32'd59606;
			5931: outdata = 32'd59605;
			5932: outdata = 32'd59604;
			5933: outdata = 32'd59603;
			5934: outdata = 32'd59602;
			5935: outdata = 32'd59601;
			5936: outdata = 32'd59600;
			5937: outdata = 32'd59599;
			5938: outdata = 32'd59598;
			5939: outdata = 32'd59597;
			5940: outdata = 32'd59596;
			5941: outdata = 32'd59595;
			5942: outdata = 32'd59594;
			5943: outdata = 32'd59593;
			5944: outdata = 32'd59592;
			5945: outdata = 32'd59591;
			5946: outdata = 32'd59590;
			5947: outdata = 32'd59589;
			5948: outdata = 32'd59588;
			5949: outdata = 32'd59587;
			5950: outdata = 32'd59586;
			5951: outdata = 32'd59585;
			5952: outdata = 32'd59584;
			5953: outdata = 32'd59583;
			5954: outdata = 32'd59582;
			5955: outdata = 32'd59581;
			5956: outdata = 32'd59580;
			5957: outdata = 32'd59579;
			5958: outdata = 32'd59578;
			5959: outdata = 32'd59577;
			5960: outdata = 32'd59576;
			5961: outdata = 32'd59575;
			5962: outdata = 32'd59574;
			5963: outdata = 32'd59573;
			5964: outdata = 32'd59572;
			5965: outdata = 32'd59571;
			5966: outdata = 32'd59570;
			5967: outdata = 32'd59569;
			5968: outdata = 32'd59568;
			5969: outdata = 32'd59567;
			5970: outdata = 32'd59566;
			5971: outdata = 32'd59565;
			5972: outdata = 32'd59564;
			5973: outdata = 32'd59563;
			5974: outdata = 32'd59562;
			5975: outdata = 32'd59561;
			5976: outdata = 32'd59560;
			5977: outdata = 32'd59559;
			5978: outdata = 32'd59558;
			5979: outdata = 32'd59557;
			5980: outdata = 32'd59556;
			5981: outdata = 32'd59555;
			5982: outdata = 32'd59554;
			5983: outdata = 32'd59553;
			5984: outdata = 32'd59552;
			5985: outdata = 32'd59551;
			5986: outdata = 32'd59550;
			5987: outdata = 32'd59549;
			5988: outdata = 32'd59548;
			5989: outdata = 32'd59547;
			5990: outdata = 32'd59546;
			5991: outdata = 32'd59545;
			5992: outdata = 32'd59544;
			5993: outdata = 32'd59543;
			5994: outdata = 32'd59542;
			5995: outdata = 32'd59541;
			5996: outdata = 32'd59540;
			5997: outdata = 32'd59539;
			5998: outdata = 32'd59538;
			5999: outdata = 32'd59537;
			6000: outdata = 32'd59536;
			6001: outdata = 32'd59535;
			6002: outdata = 32'd59534;
			6003: outdata = 32'd59533;
			6004: outdata = 32'd59532;
			6005: outdata = 32'd59531;
			6006: outdata = 32'd59530;
			6007: outdata = 32'd59529;
			6008: outdata = 32'd59528;
			6009: outdata = 32'd59527;
			6010: outdata = 32'd59526;
			6011: outdata = 32'd59525;
			6012: outdata = 32'd59524;
			6013: outdata = 32'd59523;
			6014: outdata = 32'd59522;
			6015: outdata = 32'd59521;
			6016: outdata = 32'd59520;
			6017: outdata = 32'd59519;
			6018: outdata = 32'd59518;
			6019: outdata = 32'd59517;
			6020: outdata = 32'd59516;
			6021: outdata = 32'd59515;
			6022: outdata = 32'd59514;
			6023: outdata = 32'd59513;
			6024: outdata = 32'd59512;
			6025: outdata = 32'd59511;
			6026: outdata = 32'd59510;
			6027: outdata = 32'd59509;
			6028: outdata = 32'd59508;
			6029: outdata = 32'd59507;
			6030: outdata = 32'd59506;
			6031: outdata = 32'd59505;
			6032: outdata = 32'd59504;
			6033: outdata = 32'd59503;
			6034: outdata = 32'd59502;
			6035: outdata = 32'd59501;
			6036: outdata = 32'd59500;
			6037: outdata = 32'd59499;
			6038: outdata = 32'd59498;
			6039: outdata = 32'd59497;
			6040: outdata = 32'd59496;
			6041: outdata = 32'd59495;
			6042: outdata = 32'd59494;
			6043: outdata = 32'd59493;
			6044: outdata = 32'd59492;
			6045: outdata = 32'd59491;
			6046: outdata = 32'd59490;
			6047: outdata = 32'd59489;
			6048: outdata = 32'd59488;
			6049: outdata = 32'd59487;
			6050: outdata = 32'd59486;
			6051: outdata = 32'd59485;
			6052: outdata = 32'd59484;
			6053: outdata = 32'd59483;
			6054: outdata = 32'd59482;
			6055: outdata = 32'd59481;
			6056: outdata = 32'd59480;
			6057: outdata = 32'd59479;
			6058: outdata = 32'd59478;
			6059: outdata = 32'd59477;
			6060: outdata = 32'd59476;
			6061: outdata = 32'd59475;
			6062: outdata = 32'd59474;
			6063: outdata = 32'd59473;
			6064: outdata = 32'd59472;
			6065: outdata = 32'd59471;
			6066: outdata = 32'd59470;
			6067: outdata = 32'd59469;
			6068: outdata = 32'd59468;
			6069: outdata = 32'd59467;
			6070: outdata = 32'd59466;
			6071: outdata = 32'd59465;
			6072: outdata = 32'd59464;
			6073: outdata = 32'd59463;
			6074: outdata = 32'd59462;
			6075: outdata = 32'd59461;
			6076: outdata = 32'd59460;
			6077: outdata = 32'd59459;
			6078: outdata = 32'd59458;
			6079: outdata = 32'd59457;
			6080: outdata = 32'd59456;
			6081: outdata = 32'd59455;
			6082: outdata = 32'd59454;
			6083: outdata = 32'd59453;
			6084: outdata = 32'd59452;
			6085: outdata = 32'd59451;
			6086: outdata = 32'd59450;
			6087: outdata = 32'd59449;
			6088: outdata = 32'd59448;
			6089: outdata = 32'd59447;
			6090: outdata = 32'd59446;
			6091: outdata = 32'd59445;
			6092: outdata = 32'd59444;
			6093: outdata = 32'd59443;
			6094: outdata = 32'd59442;
			6095: outdata = 32'd59441;
			6096: outdata = 32'd59440;
			6097: outdata = 32'd59439;
			6098: outdata = 32'd59438;
			6099: outdata = 32'd59437;
			6100: outdata = 32'd59436;
			6101: outdata = 32'd59435;
			6102: outdata = 32'd59434;
			6103: outdata = 32'd59433;
			6104: outdata = 32'd59432;
			6105: outdata = 32'd59431;
			6106: outdata = 32'd59430;
			6107: outdata = 32'd59429;
			6108: outdata = 32'd59428;
			6109: outdata = 32'd59427;
			6110: outdata = 32'd59426;
			6111: outdata = 32'd59425;
			6112: outdata = 32'd59424;
			6113: outdata = 32'd59423;
			6114: outdata = 32'd59422;
			6115: outdata = 32'd59421;
			6116: outdata = 32'd59420;
			6117: outdata = 32'd59419;
			6118: outdata = 32'd59418;
			6119: outdata = 32'd59417;
			6120: outdata = 32'd59416;
			6121: outdata = 32'd59415;
			6122: outdata = 32'd59414;
			6123: outdata = 32'd59413;
			6124: outdata = 32'd59412;
			6125: outdata = 32'd59411;
			6126: outdata = 32'd59410;
			6127: outdata = 32'd59409;
			6128: outdata = 32'd59408;
			6129: outdata = 32'd59407;
			6130: outdata = 32'd59406;
			6131: outdata = 32'd59405;
			6132: outdata = 32'd59404;
			6133: outdata = 32'd59403;
			6134: outdata = 32'd59402;
			6135: outdata = 32'd59401;
			6136: outdata = 32'd59400;
			6137: outdata = 32'd59399;
			6138: outdata = 32'd59398;
			6139: outdata = 32'd59397;
			6140: outdata = 32'd59396;
			6141: outdata = 32'd59395;
			6142: outdata = 32'd59394;
			6143: outdata = 32'd59393;
			6144: outdata = 32'd59392;
			6145: outdata = 32'd59391;
			6146: outdata = 32'd59390;
			6147: outdata = 32'd59389;
			6148: outdata = 32'd59388;
			6149: outdata = 32'd59387;
			6150: outdata = 32'd59386;
			6151: outdata = 32'd59385;
			6152: outdata = 32'd59384;
			6153: outdata = 32'd59383;
			6154: outdata = 32'd59382;
			6155: outdata = 32'd59381;
			6156: outdata = 32'd59380;
			6157: outdata = 32'd59379;
			6158: outdata = 32'd59378;
			6159: outdata = 32'd59377;
			6160: outdata = 32'd59376;
			6161: outdata = 32'd59375;
			6162: outdata = 32'd59374;
			6163: outdata = 32'd59373;
			6164: outdata = 32'd59372;
			6165: outdata = 32'd59371;
			6166: outdata = 32'd59370;
			6167: outdata = 32'd59369;
			6168: outdata = 32'd59368;
			6169: outdata = 32'd59367;
			6170: outdata = 32'd59366;
			6171: outdata = 32'd59365;
			6172: outdata = 32'd59364;
			6173: outdata = 32'd59363;
			6174: outdata = 32'd59362;
			6175: outdata = 32'd59361;
			6176: outdata = 32'd59360;
			6177: outdata = 32'd59359;
			6178: outdata = 32'd59358;
			6179: outdata = 32'd59357;
			6180: outdata = 32'd59356;
			6181: outdata = 32'd59355;
			6182: outdata = 32'd59354;
			6183: outdata = 32'd59353;
			6184: outdata = 32'd59352;
			6185: outdata = 32'd59351;
			6186: outdata = 32'd59350;
			6187: outdata = 32'd59349;
			6188: outdata = 32'd59348;
			6189: outdata = 32'd59347;
			6190: outdata = 32'd59346;
			6191: outdata = 32'd59345;
			6192: outdata = 32'd59344;
			6193: outdata = 32'd59343;
			6194: outdata = 32'd59342;
			6195: outdata = 32'd59341;
			6196: outdata = 32'd59340;
			6197: outdata = 32'd59339;
			6198: outdata = 32'd59338;
			6199: outdata = 32'd59337;
			6200: outdata = 32'd59336;
			6201: outdata = 32'd59335;
			6202: outdata = 32'd59334;
			6203: outdata = 32'd59333;
			6204: outdata = 32'd59332;
			6205: outdata = 32'd59331;
			6206: outdata = 32'd59330;
			6207: outdata = 32'd59329;
			6208: outdata = 32'd59328;
			6209: outdata = 32'd59327;
			6210: outdata = 32'd59326;
			6211: outdata = 32'd59325;
			6212: outdata = 32'd59324;
			6213: outdata = 32'd59323;
			6214: outdata = 32'd59322;
			6215: outdata = 32'd59321;
			6216: outdata = 32'd59320;
			6217: outdata = 32'd59319;
			6218: outdata = 32'd59318;
			6219: outdata = 32'd59317;
			6220: outdata = 32'd59316;
			6221: outdata = 32'd59315;
			6222: outdata = 32'd59314;
			6223: outdata = 32'd59313;
			6224: outdata = 32'd59312;
			6225: outdata = 32'd59311;
			6226: outdata = 32'd59310;
			6227: outdata = 32'd59309;
			6228: outdata = 32'd59308;
			6229: outdata = 32'd59307;
			6230: outdata = 32'd59306;
			6231: outdata = 32'd59305;
			6232: outdata = 32'd59304;
			6233: outdata = 32'd59303;
			6234: outdata = 32'd59302;
			6235: outdata = 32'd59301;
			6236: outdata = 32'd59300;
			6237: outdata = 32'd59299;
			6238: outdata = 32'd59298;
			6239: outdata = 32'd59297;
			6240: outdata = 32'd59296;
			6241: outdata = 32'd59295;
			6242: outdata = 32'd59294;
			6243: outdata = 32'd59293;
			6244: outdata = 32'd59292;
			6245: outdata = 32'd59291;
			6246: outdata = 32'd59290;
			6247: outdata = 32'd59289;
			6248: outdata = 32'd59288;
			6249: outdata = 32'd59287;
			6250: outdata = 32'd59286;
			6251: outdata = 32'd59285;
			6252: outdata = 32'd59284;
			6253: outdata = 32'd59283;
			6254: outdata = 32'd59282;
			6255: outdata = 32'd59281;
			6256: outdata = 32'd59280;
			6257: outdata = 32'd59279;
			6258: outdata = 32'd59278;
			6259: outdata = 32'd59277;
			6260: outdata = 32'd59276;
			6261: outdata = 32'd59275;
			6262: outdata = 32'd59274;
			6263: outdata = 32'd59273;
			6264: outdata = 32'd59272;
			6265: outdata = 32'd59271;
			6266: outdata = 32'd59270;
			6267: outdata = 32'd59269;
			6268: outdata = 32'd59268;
			6269: outdata = 32'd59267;
			6270: outdata = 32'd59266;
			6271: outdata = 32'd59265;
			6272: outdata = 32'd59264;
			6273: outdata = 32'd59263;
			6274: outdata = 32'd59262;
			6275: outdata = 32'd59261;
			6276: outdata = 32'd59260;
			6277: outdata = 32'd59259;
			6278: outdata = 32'd59258;
			6279: outdata = 32'd59257;
			6280: outdata = 32'd59256;
			6281: outdata = 32'd59255;
			6282: outdata = 32'd59254;
			6283: outdata = 32'd59253;
			6284: outdata = 32'd59252;
			6285: outdata = 32'd59251;
			6286: outdata = 32'd59250;
			6287: outdata = 32'd59249;
			6288: outdata = 32'd59248;
			6289: outdata = 32'd59247;
			6290: outdata = 32'd59246;
			6291: outdata = 32'd59245;
			6292: outdata = 32'd59244;
			6293: outdata = 32'd59243;
			6294: outdata = 32'd59242;
			6295: outdata = 32'd59241;
			6296: outdata = 32'd59240;
			6297: outdata = 32'd59239;
			6298: outdata = 32'd59238;
			6299: outdata = 32'd59237;
			6300: outdata = 32'd59236;
			6301: outdata = 32'd59235;
			6302: outdata = 32'd59234;
			6303: outdata = 32'd59233;
			6304: outdata = 32'd59232;
			6305: outdata = 32'd59231;
			6306: outdata = 32'd59230;
			6307: outdata = 32'd59229;
			6308: outdata = 32'd59228;
			6309: outdata = 32'd59227;
			6310: outdata = 32'd59226;
			6311: outdata = 32'd59225;
			6312: outdata = 32'd59224;
			6313: outdata = 32'd59223;
			6314: outdata = 32'd59222;
			6315: outdata = 32'd59221;
			6316: outdata = 32'd59220;
			6317: outdata = 32'd59219;
			6318: outdata = 32'd59218;
			6319: outdata = 32'd59217;
			6320: outdata = 32'd59216;
			6321: outdata = 32'd59215;
			6322: outdata = 32'd59214;
			6323: outdata = 32'd59213;
			6324: outdata = 32'd59212;
			6325: outdata = 32'd59211;
			6326: outdata = 32'd59210;
			6327: outdata = 32'd59209;
			6328: outdata = 32'd59208;
			6329: outdata = 32'd59207;
			6330: outdata = 32'd59206;
			6331: outdata = 32'd59205;
			6332: outdata = 32'd59204;
			6333: outdata = 32'd59203;
			6334: outdata = 32'd59202;
			6335: outdata = 32'd59201;
			6336: outdata = 32'd59200;
			6337: outdata = 32'd59199;
			6338: outdata = 32'd59198;
			6339: outdata = 32'd59197;
			6340: outdata = 32'd59196;
			6341: outdata = 32'd59195;
			6342: outdata = 32'd59194;
			6343: outdata = 32'd59193;
			6344: outdata = 32'd59192;
			6345: outdata = 32'd59191;
			6346: outdata = 32'd59190;
			6347: outdata = 32'd59189;
			6348: outdata = 32'd59188;
			6349: outdata = 32'd59187;
			6350: outdata = 32'd59186;
			6351: outdata = 32'd59185;
			6352: outdata = 32'd59184;
			6353: outdata = 32'd59183;
			6354: outdata = 32'd59182;
			6355: outdata = 32'd59181;
			6356: outdata = 32'd59180;
			6357: outdata = 32'd59179;
			6358: outdata = 32'd59178;
			6359: outdata = 32'd59177;
			6360: outdata = 32'd59176;
			6361: outdata = 32'd59175;
			6362: outdata = 32'd59174;
			6363: outdata = 32'd59173;
			6364: outdata = 32'd59172;
			6365: outdata = 32'd59171;
			6366: outdata = 32'd59170;
			6367: outdata = 32'd59169;
			6368: outdata = 32'd59168;
			6369: outdata = 32'd59167;
			6370: outdata = 32'd59166;
			6371: outdata = 32'd59165;
			6372: outdata = 32'd59164;
			6373: outdata = 32'd59163;
			6374: outdata = 32'd59162;
			6375: outdata = 32'd59161;
			6376: outdata = 32'd59160;
			6377: outdata = 32'd59159;
			6378: outdata = 32'd59158;
			6379: outdata = 32'd59157;
			6380: outdata = 32'd59156;
			6381: outdata = 32'd59155;
			6382: outdata = 32'd59154;
			6383: outdata = 32'd59153;
			6384: outdata = 32'd59152;
			6385: outdata = 32'd59151;
			6386: outdata = 32'd59150;
			6387: outdata = 32'd59149;
			6388: outdata = 32'd59148;
			6389: outdata = 32'd59147;
			6390: outdata = 32'd59146;
			6391: outdata = 32'd59145;
			6392: outdata = 32'd59144;
			6393: outdata = 32'd59143;
			6394: outdata = 32'd59142;
			6395: outdata = 32'd59141;
			6396: outdata = 32'd59140;
			6397: outdata = 32'd59139;
			6398: outdata = 32'd59138;
			6399: outdata = 32'd59137;
			6400: outdata = 32'd59136;
			6401: outdata = 32'd59135;
			6402: outdata = 32'd59134;
			6403: outdata = 32'd59133;
			6404: outdata = 32'd59132;
			6405: outdata = 32'd59131;
			6406: outdata = 32'd59130;
			6407: outdata = 32'd59129;
			6408: outdata = 32'd59128;
			6409: outdata = 32'd59127;
			6410: outdata = 32'd59126;
			6411: outdata = 32'd59125;
			6412: outdata = 32'd59124;
			6413: outdata = 32'd59123;
			6414: outdata = 32'd59122;
			6415: outdata = 32'd59121;
			6416: outdata = 32'd59120;
			6417: outdata = 32'd59119;
			6418: outdata = 32'd59118;
			6419: outdata = 32'd59117;
			6420: outdata = 32'd59116;
			6421: outdata = 32'd59115;
			6422: outdata = 32'd59114;
			6423: outdata = 32'd59113;
			6424: outdata = 32'd59112;
			6425: outdata = 32'd59111;
			6426: outdata = 32'd59110;
			6427: outdata = 32'd59109;
			6428: outdata = 32'd59108;
			6429: outdata = 32'd59107;
			6430: outdata = 32'd59106;
			6431: outdata = 32'd59105;
			6432: outdata = 32'd59104;
			6433: outdata = 32'd59103;
			6434: outdata = 32'd59102;
			6435: outdata = 32'd59101;
			6436: outdata = 32'd59100;
			6437: outdata = 32'd59099;
			6438: outdata = 32'd59098;
			6439: outdata = 32'd59097;
			6440: outdata = 32'd59096;
			6441: outdata = 32'd59095;
			6442: outdata = 32'd59094;
			6443: outdata = 32'd59093;
			6444: outdata = 32'd59092;
			6445: outdata = 32'd59091;
			6446: outdata = 32'd59090;
			6447: outdata = 32'd59089;
			6448: outdata = 32'd59088;
			6449: outdata = 32'd59087;
			6450: outdata = 32'd59086;
			6451: outdata = 32'd59085;
			6452: outdata = 32'd59084;
			6453: outdata = 32'd59083;
			6454: outdata = 32'd59082;
			6455: outdata = 32'd59081;
			6456: outdata = 32'd59080;
			6457: outdata = 32'd59079;
			6458: outdata = 32'd59078;
			6459: outdata = 32'd59077;
			6460: outdata = 32'd59076;
			6461: outdata = 32'd59075;
			6462: outdata = 32'd59074;
			6463: outdata = 32'd59073;
			6464: outdata = 32'd59072;
			6465: outdata = 32'd59071;
			6466: outdata = 32'd59070;
			6467: outdata = 32'd59069;
			6468: outdata = 32'd59068;
			6469: outdata = 32'd59067;
			6470: outdata = 32'd59066;
			6471: outdata = 32'd59065;
			6472: outdata = 32'd59064;
			6473: outdata = 32'd59063;
			6474: outdata = 32'd59062;
			6475: outdata = 32'd59061;
			6476: outdata = 32'd59060;
			6477: outdata = 32'd59059;
			6478: outdata = 32'd59058;
			6479: outdata = 32'd59057;
			6480: outdata = 32'd59056;
			6481: outdata = 32'd59055;
			6482: outdata = 32'd59054;
			6483: outdata = 32'd59053;
			6484: outdata = 32'd59052;
			6485: outdata = 32'd59051;
			6486: outdata = 32'd59050;
			6487: outdata = 32'd59049;
			6488: outdata = 32'd59048;
			6489: outdata = 32'd59047;
			6490: outdata = 32'd59046;
			6491: outdata = 32'd59045;
			6492: outdata = 32'd59044;
			6493: outdata = 32'd59043;
			6494: outdata = 32'd59042;
			6495: outdata = 32'd59041;
			6496: outdata = 32'd59040;
			6497: outdata = 32'd59039;
			6498: outdata = 32'd59038;
			6499: outdata = 32'd59037;
			6500: outdata = 32'd59036;
			6501: outdata = 32'd59035;
			6502: outdata = 32'd59034;
			6503: outdata = 32'd59033;
			6504: outdata = 32'd59032;
			6505: outdata = 32'd59031;
			6506: outdata = 32'd59030;
			6507: outdata = 32'd59029;
			6508: outdata = 32'd59028;
			6509: outdata = 32'd59027;
			6510: outdata = 32'd59026;
			6511: outdata = 32'd59025;
			6512: outdata = 32'd59024;
			6513: outdata = 32'd59023;
			6514: outdata = 32'd59022;
			6515: outdata = 32'd59021;
			6516: outdata = 32'd59020;
			6517: outdata = 32'd59019;
			6518: outdata = 32'd59018;
			6519: outdata = 32'd59017;
			6520: outdata = 32'd59016;
			6521: outdata = 32'd59015;
			6522: outdata = 32'd59014;
			6523: outdata = 32'd59013;
			6524: outdata = 32'd59012;
			6525: outdata = 32'd59011;
			6526: outdata = 32'd59010;
			6527: outdata = 32'd59009;
			6528: outdata = 32'd59008;
			6529: outdata = 32'd59007;
			6530: outdata = 32'd59006;
			6531: outdata = 32'd59005;
			6532: outdata = 32'd59004;
			6533: outdata = 32'd59003;
			6534: outdata = 32'd59002;
			6535: outdata = 32'd59001;
			6536: outdata = 32'd59000;
			6537: outdata = 32'd58999;
			6538: outdata = 32'd58998;
			6539: outdata = 32'd58997;
			6540: outdata = 32'd58996;
			6541: outdata = 32'd58995;
			6542: outdata = 32'd58994;
			6543: outdata = 32'd58993;
			6544: outdata = 32'd58992;
			6545: outdata = 32'd58991;
			6546: outdata = 32'd58990;
			6547: outdata = 32'd58989;
			6548: outdata = 32'd58988;
			6549: outdata = 32'd58987;
			6550: outdata = 32'd58986;
			6551: outdata = 32'd58985;
			6552: outdata = 32'd58984;
			6553: outdata = 32'd58983;
			6554: outdata = 32'd58982;
			6555: outdata = 32'd58981;
			6556: outdata = 32'd58980;
			6557: outdata = 32'd58979;
			6558: outdata = 32'd58978;
			6559: outdata = 32'd58977;
			6560: outdata = 32'd58976;
			6561: outdata = 32'd58975;
			6562: outdata = 32'd58974;
			6563: outdata = 32'd58973;
			6564: outdata = 32'd58972;
			6565: outdata = 32'd58971;
			6566: outdata = 32'd58970;
			6567: outdata = 32'd58969;
			6568: outdata = 32'd58968;
			6569: outdata = 32'd58967;
			6570: outdata = 32'd58966;
			6571: outdata = 32'd58965;
			6572: outdata = 32'd58964;
			6573: outdata = 32'd58963;
			6574: outdata = 32'd58962;
			6575: outdata = 32'd58961;
			6576: outdata = 32'd58960;
			6577: outdata = 32'd58959;
			6578: outdata = 32'd58958;
			6579: outdata = 32'd58957;
			6580: outdata = 32'd58956;
			6581: outdata = 32'd58955;
			6582: outdata = 32'd58954;
			6583: outdata = 32'd58953;
			6584: outdata = 32'd58952;
			6585: outdata = 32'd58951;
			6586: outdata = 32'd58950;
			6587: outdata = 32'd58949;
			6588: outdata = 32'd58948;
			6589: outdata = 32'd58947;
			6590: outdata = 32'd58946;
			6591: outdata = 32'd58945;
			6592: outdata = 32'd58944;
			6593: outdata = 32'd58943;
			6594: outdata = 32'd58942;
			6595: outdata = 32'd58941;
			6596: outdata = 32'd58940;
			6597: outdata = 32'd58939;
			6598: outdata = 32'd58938;
			6599: outdata = 32'd58937;
			6600: outdata = 32'd58936;
			6601: outdata = 32'd58935;
			6602: outdata = 32'd58934;
			6603: outdata = 32'd58933;
			6604: outdata = 32'd58932;
			6605: outdata = 32'd58931;
			6606: outdata = 32'd58930;
			6607: outdata = 32'd58929;
			6608: outdata = 32'd58928;
			6609: outdata = 32'd58927;
			6610: outdata = 32'd58926;
			6611: outdata = 32'd58925;
			6612: outdata = 32'd58924;
			6613: outdata = 32'd58923;
			6614: outdata = 32'd58922;
			6615: outdata = 32'd58921;
			6616: outdata = 32'd58920;
			6617: outdata = 32'd58919;
			6618: outdata = 32'd58918;
			6619: outdata = 32'd58917;
			6620: outdata = 32'd58916;
			6621: outdata = 32'd58915;
			6622: outdata = 32'd58914;
			6623: outdata = 32'd58913;
			6624: outdata = 32'd58912;
			6625: outdata = 32'd58911;
			6626: outdata = 32'd58910;
			6627: outdata = 32'd58909;
			6628: outdata = 32'd58908;
			6629: outdata = 32'd58907;
			6630: outdata = 32'd58906;
			6631: outdata = 32'd58905;
			6632: outdata = 32'd58904;
			6633: outdata = 32'd58903;
			6634: outdata = 32'd58902;
			6635: outdata = 32'd58901;
			6636: outdata = 32'd58900;
			6637: outdata = 32'd58899;
			6638: outdata = 32'd58898;
			6639: outdata = 32'd58897;
			6640: outdata = 32'd58896;
			6641: outdata = 32'd58895;
			6642: outdata = 32'd58894;
			6643: outdata = 32'd58893;
			6644: outdata = 32'd58892;
			6645: outdata = 32'd58891;
			6646: outdata = 32'd58890;
			6647: outdata = 32'd58889;
			6648: outdata = 32'd58888;
			6649: outdata = 32'd58887;
			6650: outdata = 32'd58886;
			6651: outdata = 32'd58885;
			6652: outdata = 32'd58884;
			6653: outdata = 32'd58883;
			6654: outdata = 32'd58882;
			6655: outdata = 32'd58881;
			6656: outdata = 32'd58880;
			6657: outdata = 32'd58879;
			6658: outdata = 32'd58878;
			6659: outdata = 32'd58877;
			6660: outdata = 32'd58876;
			6661: outdata = 32'd58875;
			6662: outdata = 32'd58874;
			6663: outdata = 32'd58873;
			6664: outdata = 32'd58872;
			6665: outdata = 32'd58871;
			6666: outdata = 32'd58870;
			6667: outdata = 32'd58869;
			6668: outdata = 32'd58868;
			6669: outdata = 32'd58867;
			6670: outdata = 32'd58866;
			6671: outdata = 32'd58865;
			6672: outdata = 32'd58864;
			6673: outdata = 32'd58863;
			6674: outdata = 32'd58862;
			6675: outdata = 32'd58861;
			6676: outdata = 32'd58860;
			6677: outdata = 32'd58859;
			6678: outdata = 32'd58858;
			6679: outdata = 32'd58857;
			6680: outdata = 32'd58856;
			6681: outdata = 32'd58855;
			6682: outdata = 32'd58854;
			6683: outdata = 32'd58853;
			6684: outdata = 32'd58852;
			6685: outdata = 32'd58851;
			6686: outdata = 32'd58850;
			6687: outdata = 32'd58849;
			6688: outdata = 32'd58848;
			6689: outdata = 32'd58847;
			6690: outdata = 32'd58846;
			6691: outdata = 32'd58845;
			6692: outdata = 32'd58844;
			6693: outdata = 32'd58843;
			6694: outdata = 32'd58842;
			6695: outdata = 32'd58841;
			6696: outdata = 32'd58840;
			6697: outdata = 32'd58839;
			6698: outdata = 32'd58838;
			6699: outdata = 32'd58837;
			6700: outdata = 32'd58836;
			6701: outdata = 32'd58835;
			6702: outdata = 32'd58834;
			6703: outdata = 32'd58833;
			6704: outdata = 32'd58832;
			6705: outdata = 32'd58831;
			6706: outdata = 32'd58830;
			6707: outdata = 32'd58829;
			6708: outdata = 32'd58828;
			6709: outdata = 32'd58827;
			6710: outdata = 32'd58826;
			6711: outdata = 32'd58825;
			6712: outdata = 32'd58824;
			6713: outdata = 32'd58823;
			6714: outdata = 32'd58822;
			6715: outdata = 32'd58821;
			6716: outdata = 32'd58820;
			6717: outdata = 32'd58819;
			6718: outdata = 32'd58818;
			6719: outdata = 32'd58817;
			6720: outdata = 32'd58816;
			6721: outdata = 32'd58815;
			6722: outdata = 32'd58814;
			6723: outdata = 32'd58813;
			6724: outdata = 32'd58812;
			6725: outdata = 32'd58811;
			6726: outdata = 32'd58810;
			6727: outdata = 32'd58809;
			6728: outdata = 32'd58808;
			6729: outdata = 32'd58807;
			6730: outdata = 32'd58806;
			6731: outdata = 32'd58805;
			6732: outdata = 32'd58804;
			6733: outdata = 32'd58803;
			6734: outdata = 32'd58802;
			6735: outdata = 32'd58801;
			6736: outdata = 32'd58800;
			6737: outdata = 32'd58799;
			6738: outdata = 32'd58798;
			6739: outdata = 32'd58797;
			6740: outdata = 32'd58796;
			6741: outdata = 32'd58795;
			6742: outdata = 32'd58794;
			6743: outdata = 32'd58793;
			6744: outdata = 32'd58792;
			6745: outdata = 32'd58791;
			6746: outdata = 32'd58790;
			6747: outdata = 32'd58789;
			6748: outdata = 32'd58788;
			6749: outdata = 32'd58787;
			6750: outdata = 32'd58786;
			6751: outdata = 32'd58785;
			6752: outdata = 32'd58784;
			6753: outdata = 32'd58783;
			6754: outdata = 32'd58782;
			6755: outdata = 32'd58781;
			6756: outdata = 32'd58780;
			6757: outdata = 32'd58779;
			6758: outdata = 32'd58778;
			6759: outdata = 32'd58777;
			6760: outdata = 32'd58776;
			6761: outdata = 32'd58775;
			6762: outdata = 32'd58774;
			6763: outdata = 32'd58773;
			6764: outdata = 32'd58772;
			6765: outdata = 32'd58771;
			6766: outdata = 32'd58770;
			6767: outdata = 32'd58769;
			6768: outdata = 32'd58768;
			6769: outdata = 32'd58767;
			6770: outdata = 32'd58766;
			6771: outdata = 32'd58765;
			6772: outdata = 32'd58764;
			6773: outdata = 32'd58763;
			6774: outdata = 32'd58762;
			6775: outdata = 32'd58761;
			6776: outdata = 32'd58760;
			6777: outdata = 32'd58759;
			6778: outdata = 32'd58758;
			6779: outdata = 32'd58757;
			6780: outdata = 32'd58756;
			6781: outdata = 32'd58755;
			6782: outdata = 32'd58754;
			6783: outdata = 32'd58753;
			6784: outdata = 32'd58752;
			6785: outdata = 32'd58751;
			6786: outdata = 32'd58750;
			6787: outdata = 32'd58749;
			6788: outdata = 32'd58748;
			6789: outdata = 32'd58747;
			6790: outdata = 32'd58746;
			6791: outdata = 32'd58745;
			6792: outdata = 32'd58744;
			6793: outdata = 32'd58743;
			6794: outdata = 32'd58742;
			6795: outdata = 32'd58741;
			6796: outdata = 32'd58740;
			6797: outdata = 32'd58739;
			6798: outdata = 32'd58738;
			6799: outdata = 32'd58737;
			6800: outdata = 32'd58736;
			6801: outdata = 32'd58735;
			6802: outdata = 32'd58734;
			6803: outdata = 32'd58733;
			6804: outdata = 32'd58732;
			6805: outdata = 32'd58731;
			6806: outdata = 32'd58730;
			6807: outdata = 32'd58729;
			6808: outdata = 32'd58728;
			6809: outdata = 32'd58727;
			6810: outdata = 32'd58726;
			6811: outdata = 32'd58725;
			6812: outdata = 32'd58724;
			6813: outdata = 32'd58723;
			6814: outdata = 32'd58722;
			6815: outdata = 32'd58721;
			6816: outdata = 32'd58720;
			6817: outdata = 32'd58719;
			6818: outdata = 32'd58718;
			6819: outdata = 32'd58717;
			6820: outdata = 32'd58716;
			6821: outdata = 32'd58715;
			6822: outdata = 32'd58714;
			6823: outdata = 32'd58713;
			6824: outdata = 32'd58712;
			6825: outdata = 32'd58711;
			6826: outdata = 32'd58710;
			6827: outdata = 32'd58709;
			6828: outdata = 32'd58708;
			6829: outdata = 32'd58707;
			6830: outdata = 32'd58706;
			6831: outdata = 32'd58705;
			6832: outdata = 32'd58704;
			6833: outdata = 32'd58703;
			6834: outdata = 32'd58702;
			6835: outdata = 32'd58701;
			6836: outdata = 32'd58700;
			6837: outdata = 32'd58699;
			6838: outdata = 32'd58698;
			6839: outdata = 32'd58697;
			6840: outdata = 32'd58696;
			6841: outdata = 32'd58695;
			6842: outdata = 32'd58694;
			6843: outdata = 32'd58693;
			6844: outdata = 32'd58692;
			6845: outdata = 32'd58691;
			6846: outdata = 32'd58690;
			6847: outdata = 32'd58689;
			6848: outdata = 32'd58688;
			6849: outdata = 32'd58687;
			6850: outdata = 32'd58686;
			6851: outdata = 32'd58685;
			6852: outdata = 32'd58684;
			6853: outdata = 32'd58683;
			6854: outdata = 32'd58682;
			6855: outdata = 32'd58681;
			6856: outdata = 32'd58680;
			6857: outdata = 32'd58679;
			6858: outdata = 32'd58678;
			6859: outdata = 32'd58677;
			6860: outdata = 32'd58676;
			6861: outdata = 32'd58675;
			6862: outdata = 32'd58674;
			6863: outdata = 32'd58673;
			6864: outdata = 32'd58672;
			6865: outdata = 32'd58671;
			6866: outdata = 32'd58670;
			6867: outdata = 32'd58669;
			6868: outdata = 32'd58668;
			6869: outdata = 32'd58667;
			6870: outdata = 32'd58666;
			6871: outdata = 32'd58665;
			6872: outdata = 32'd58664;
			6873: outdata = 32'd58663;
			6874: outdata = 32'd58662;
			6875: outdata = 32'd58661;
			6876: outdata = 32'd58660;
			6877: outdata = 32'd58659;
			6878: outdata = 32'd58658;
			6879: outdata = 32'd58657;
			6880: outdata = 32'd58656;
			6881: outdata = 32'd58655;
			6882: outdata = 32'd58654;
			6883: outdata = 32'd58653;
			6884: outdata = 32'd58652;
			6885: outdata = 32'd58651;
			6886: outdata = 32'd58650;
			6887: outdata = 32'd58649;
			6888: outdata = 32'd58648;
			6889: outdata = 32'd58647;
			6890: outdata = 32'd58646;
			6891: outdata = 32'd58645;
			6892: outdata = 32'd58644;
			6893: outdata = 32'd58643;
			6894: outdata = 32'd58642;
			6895: outdata = 32'd58641;
			6896: outdata = 32'd58640;
			6897: outdata = 32'd58639;
			6898: outdata = 32'd58638;
			6899: outdata = 32'd58637;
			6900: outdata = 32'd58636;
			6901: outdata = 32'd58635;
			6902: outdata = 32'd58634;
			6903: outdata = 32'd58633;
			6904: outdata = 32'd58632;
			6905: outdata = 32'd58631;
			6906: outdata = 32'd58630;
			6907: outdata = 32'd58629;
			6908: outdata = 32'd58628;
			6909: outdata = 32'd58627;
			6910: outdata = 32'd58626;
			6911: outdata = 32'd58625;
			6912: outdata = 32'd58624;
			6913: outdata = 32'd58623;
			6914: outdata = 32'd58622;
			6915: outdata = 32'd58621;
			6916: outdata = 32'd58620;
			6917: outdata = 32'd58619;
			6918: outdata = 32'd58618;
			6919: outdata = 32'd58617;
			6920: outdata = 32'd58616;
			6921: outdata = 32'd58615;
			6922: outdata = 32'd58614;
			6923: outdata = 32'd58613;
			6924: outdata = 32'd58612;
			6925: outdata = 32'd58611;
			6926: outdata = 32'd58610;
			6927: outdata = 32'd58609;
			6928: outdata = 32'd58608;
			6929: outdata = 32'd58607;
			6930: outdata = 32'd58606;
			6931: outdata = 32'd58605;
			6932: outdata = 32'd58604;
			6933: outdata = 32'd58603;
			6934: outdata = 32'd58602;
			6935: outdata = 32'd58601;
			6936: outdata = 32'd58600;
			6937: outdata = 32'd58599;
			6938: outdata = 32'd58598;
			6939: outdata = 32'd58597;
			6940: outdata = 32'd58596;
			6941: outdata = 32'd58595;
			6942: outdata = 32'd58594;
			6943: outdata = 32'd58593;
			6944: outdata = 32'd58592;
			6945: outdata = 32'd58591;
			6946: outdata = 32'd58590;
			6947: outdata = 32'd58589;
			6948: outdata = 32'd58588;
			6949: outdata = 32'd58587;
			6950: outdata = 32'd58586;
			6951: outdata = 32'd58585;
			6952: outdata = 32'd58584;
			6953: outdata = 32'd58583;
			6954: outdata = 32'd58582;
			6955: outdata = 32'd58581;
			6956: outdata = 32'd58580;
			6957: outdata = 32'd58579;
			6958: outdata = 32'd58578;
			6959: outdata = 32'd58577;
			6960: outdata = 32'd58576;
			6961: outdata = 32'd58575;
			6962: outdata = 32'd58574;
			6963: outdata = 32'd58573;
			6964: outdata = 32'd58572;
			6965: outdata = 32'd58571;
			6966: outdata = 32'd58570;
			6967: outdata = 32'd58569;
			6968: outdata = 32'd58568;
			6969: outdata = 32'd58567;
			6970: outdata = 32'd58566;
			6971: outdata = 32'd58565;
			6972: outdata = 32'd58564;
			6973: outdata = 32'd58563;
			6974: outdata = 32'd58562;
			6975: outdata = 32'd58561;
			6976: outdata = 32'd58560;
			6977: outdata = 32'd58559;
			6978: outdata = 32'd58558;
			6979: outdata = 32'd58557;
			6980: outdata = 32'd58556;
			6981: outdata = 32'd58555;
			6982: outdata = 32'd58554;
			6983: outdata = 32'd58553;
			6984: outdata = 32'd58552;
			6985: outdata = 32'd58551;
			6986: outdata = 32'd58550;
			6987: outdata = 32'd58549;
			6988: outdata = 32'd58548;
			6989: outdata = 32'd58547;
			6990: outdata = 32'd58546;
			6991: outdata = 32'd58545;
			6992: outdata = 32'd58544;
			6993: outdata = 32'd58543;
			6994: outdata = 32'd58542;
			6995: outdata = 32'd58541;
			6996: outdata = 32'd58540;
			6997: outdata = 32'd58539;
			6998: outdata = 32'd58538;
			6999: outdata = 32'd58537;
			7000: outdata = 32'd58536;
			7001: outdata = 32'd58535;
			7002: outdata = 32'd58534;
			7003: outdata = 32'd58533;
			7004: outdata = 32'd58532;
			7005: outdata = 32'd58531;
			7006: outdata = 32'd58530;
			7007: outdata = 32'd58529;
			7008: outdata = 32'd58528;
			7009: outdata = 32'd58527;
			7010: outdata = 32'd58526;
			7011: outdata = 32'd58525;
			7012: outdata = 32'd58524;
			7013: outdata = 32'd58523;
			7014: outdata = 32'd58522;
			7015: outdata = 32'd58521;
			7016: outdata = 32'd58520;
			7017: outdata = 32'd58519;
			7018: outdata = 32'd58518;
			7019: outdata = 32'd58517;
			7020: outdata = 32'd58516;
			7021: outdata = 32'd58515;
			7022: outdata = 32'd58514;
			7023: outdata = 32'd58513;
			7024: outdata = 32'd58512;
			7025: outdata = 32'd58511;
			7026: outdata = 32'd58510;
			7027: outdata = 32'd58509;
			7028: outdata = 32'd58508;
			7029: outdata = 32'd58507;
			7030: outdata = 32'd58506;
			7031: outdata = 32'd58505;
			7032: outdata = 32'd58504;
			7033: outdata = 32'd58503;
			7034: outdata = 32'd58502;
			7035: outdata = 32'd58501;
			7036: outdata = 32'd58500;
			7037: outdata = 32'd58499;
			7038: outdata = 32'd58498;
			7039: outdata = 32'd58497;
			7040: outdata = 32'd58496;
			7041: outdata = 32'd58495;
			7042: outdata = 32'd58494;
			7043: outdata = 32'd58493;
			7044: outdata = 32'd58492;
			7045: outdata = 32'd58491;
			7046: outdata = 32'd58490;
			7047: outdata = 32'd58489;
			7048: outdata = 32'd58488;
			7049: outdata = 32'd58487;
			7050: outdata = 32'd58486;
			7051: outdata = 32'd58485;
			7052: outdata = 32'd58484;
			7053: outdata = 32'd58483;
			7054: outdata = 32'd58482;
			7055: outdata = 32'd58481;
			7056: outdata = 32'd58480;
			7057: outdata = 32'd58479;
			7058: outdata = 32'd58478;
			7059: outdata = 32'd58477;
			7060: outdata = 32'd58476;
			7061: outdata = 32'd58475;
			7062: outdata = 32'd58474;
			7063: outdata = 32'd58473;
			7064: outdata = 32'd58472;
			7065: outdata = 32'd58471;
			7066: outdata = 32'd58470;
			7067: outdata = 32'd58469;
			7068: outdata = 32'd58468;
			7069: outdata = 32'd58467;
			7070: outdata = 32'd58466;
			7071: outdata = 32'd58465;
			7072: outdata = 32'd58464;
			7073: outdata = 32'd58463;
			7074: outdata = 32'd58462;
			7075: outdata = 32'd58461;
			7076: outdata = 32'd58460;
			7077: outdata = 32'd58459;
			7078: outdata = 32'd58458;
			7079: outdata = 32'd58457;
			7080: outdata = 32'd58456;
			7081: outdata = 32'd58455;
			7082: outdata = 32'd58454;
			7083: outdata = 32'd58453;
			7084: outdata = 32'd58452;
			7085: outdata = 32'd58451;
			7086: outdata = 32'd58450;
			7087: outdata = 32'd58449;
			7088: outdata = 32'd58448;
			7089: outdata = 32'd58447;
			7090: outdata = 32'd58446;
			7091: outdata = 32'd58445;
			7092: outdata = 32'd58444;
			7093: outdata = 32'd58443;
			7094: outdata = 32'd58442;
			7095: outdata = 32'd58441;
			7096: outdata = 32'd58440;
			7097: outdata = 32'd58439;
			7098: outdata = 32'd58438;
			7099: outdata = 32'd58437;
			7100: outdata = 32'd58436;
			7101: outdata = 32'd58435;
			7102: outdata = 32'd58434;
			7103: outdata = 32'd58433;
			7104: outdata = 32'd58432;
			7105: outdata = 32'd58431;
			7106: outdata = 32'd58430;
			7107: outdata = 32'd58429;
			7108: outdata = 32'd58428;
			7109: outdata = 32'd58427;
			7110: outdata = 32'd58426;
			7111: outdata = 32'd58425;
			7112: outdata = 32'd58424;
			7113: outdata = 32'd58423;
			7114: outdata = 32'd58422;
			7115: outdata = 32'd58421;
			7116: outdata = 32'd58420;
			7117: outdata = 32'd58419;
			7118: outdata = 32'd58418;
			7119: outdata = 32'd58417;
			7120: outdata = 32'd58416;
			7121: outdata = 32'd58415;
			7122: outdata = 32'd58414;
			7123: outdata = 32'd58413;
			7124: outdata = 32'd58412;
			7125: outdata = 32'd58411;
			7126: outdata = 32'd58410;
			7127: outdata = 32'd58409;
			7128: outdata = 32'd58408;
			7129: outdata = 32'd58407;
			7130: outdata = 32'd58406;
			7131: outdata = 32'd58405;
			7132: outdata = 32'd58404;
			7133: outdata = 32'd58403;
			7134: outdata = 32'd58402;
			7135: outdata = 32'd58401;
			7136: outdata = 32'd58400;
			7137: outdata = 32'd58399;
			7138: outdata = 32'd58398;
			7139: outdata = 32'd58397;
			7140: outdata = 32'd58396;
			7141: outdata = 32'd58395;
			7142: outdata = 32'd58394;
			7143: outdata = 32'd58393;
			7144: outdata = 32'd58392;
			7145: outdata = 32'd58391;
			7146: outdata = 32'd58390;
			7147: outdata = 32'd58389;
			7148: outdata = 32'd58388;
			7149: outdata = 32'd58387;
			7150: outdata = 32'd58386;
			7151: outdata = 32'd58385;
			7152: outdata = 32'd58384;
			7153: outdata = 32'd58383;
			7154: outdata = 32'd58382;
			7155: outdata = 32'd58381;
			7156: outdata = 32'd58380;
			7157: outdata = 32'd58379;
			7158: outdata = 32'd58378;
			7159: outdata = 32'd58377;
			7160: outdata = 32'd58376;
			7161: outdata = 32'd58375;
			7162: outdata = 32'd58374;
			7163: outdata = 32'd58373;
			7164: outdata = 32'd58372;
			7165: outdata = 32'd58371;
			7166: outdata = 32'd58370;
			7167: outdata = 32'd58369;
			7168: outdata = 32'd58368;
			7169: outdata = 32'd58367;
			7170: outdata = 32'd58366;
			7171: outdata = 32'd58365;
			7172: outdata = 32'd58364;
			7173: outdata = 32'd58363;
			7174: outdata = 32'd58362;
			7175: outdata = 32'd58361;
			7176: outdata = 32'd58360;
			7177: outdata = 32'd58359;
			7178: outdata = 32'd58358;
			7179: outdata = 32'd58357;
			7180: outdata = 32'd58356;
			7181: outdata = 32'd58355;
			7182: outdata = 32'd58354;
			7183: outdata = 32'd58353;
			7184: outdata = 32'd58352;
			7185: outdata = 32'd58351;
			7186: outdata = 32'd58350;
			7187: outdata = 32'd58349;
			7188: outdata = 32'd58348;
			7189: outdata = 32'd58347;
			7190: outdata = 32'd58346;
			7191: outdata = 32'd58345;
			7192: outdata = 32'd58344;
			7193: outdata = 32'd58343;
			7194: outdata = 32'd58342;
			7195: outdata = 32'd58341;
			7196: outdata = 32'd58340;
			7197: outdata = 32'd58339;
			7198: outdata = 32'd58338;
			7199: outdata = 32'd58337;
			7200: outdata = 32'd58336;
			7201: outdata = 32'd58335;
			7202: outdata = 32'd58334;
			7203: outdata = 32'd58333;
			7204: outdata = 32'd58332;
			7205: outdata = 32'd58331;
			7206: outdata = 32'd58330;
			7207: outdata = 32'd58329;
			7208: outdata = 32'd58328;
			7209: outdata = 32'd58327;
			7210: outdata = 32'd58326;
			7211: outdata = 32'd58325;
			7212: outdata = 32'd58324;
			7213: outdata = 32'd58323;
			7214: outdata = 32'd58322;
			7215: outdata = 32'd58321;
			7216: outdata = 32'd58320;
			7217: outdata = 32'd58319;
			7218: outdata = 32'd58318;
			7219: outdata = 32'd58317;
			7220: outdata = 32'd58316;
			7221: outdata = 32'd58315;
			7222: outdata = 32'd58314;
			7223: outdata = 32'd58313;
			7224: outdata = 32'd58312;
			7225: outdata = 32'd58311;
			7226: outdata = 32'd58310;
			7227: outdata = 32'd58309;
			7228: outdata = 32'd58308;
			7229: outdata = 32'd58307;
			7230: outdata = 32'd58306;
			7231: outdata = 32'd58305;
			7232: outdata = 32'd58304;
			7233: outdata = 32'd58303;
			7234: outdata = 32'd58302;
			7235: outdata = 32'd58301;
			7236: outdata = 32'd58300;
			7237: outdata = 32'd58299;
			7238: outdata = 32'd58298;
			7239: outdata = 32'd58297;
			7240: outdata = 32'd58296;
			7241: outdata = 32'd58295;
			7242: outdata = 32'd58294;
			7243: outdata = 32'd58293;
			7244: outdata = 32'd58292;
			7245: outdata = 32'd58291;
			7246: outdata = 32'd58290;
			7247: outdata = 32'd58289;
			7248: outdata = 32'd58288;
			7249: outdata = 32'd58287;
			7250: outdata = 32'd58286;
			7251: outdata = 32'd58285;
			7252: outdata = 32'd58284;
			7253: outdata = 32'd58283;
			7254: outdata = 32'd58282;
			7255: outdata = 32'd58281;
			7256: outdata = 32'd58280;
			7257: outdata = 32'd58279;
			7258: outdata = 32'd58278;
			7259: outdata = 32'd58277;
			7260: outdata = 32'd58276;
			7261: outdata = 32'd58275;
			7262: outdata = 32'd58274;
			7263: outdata = 32'd58273;
			7264: outdata = 32'd58272;
			7265: outdata = 32'd58271;
			7266: outdata = 32'd58270;
			7267: outdata = 32'd58269;
			7268: outdata = 32'd58268;
			7269: outdata = 32'd58267;
			7270: outdata = 32'd58266;
			7271: outdata = 32'd58265;
			7272: outdata = 32'd58264;
			7273: outdata = 32'd58263;
			7274: outdata = 32'd58262;
			7275: outdata = 32'd58261;
			7276: outdata = 32'd58260;
			7277: outdata = 32'd58259;
			7278: outdata = 32'd58258;
			7279: outdata = 32'd58257;
			7280: outdata = 32'd58256;
			7281: outdata = 32'd58255;
			7282: outdata = 32'd58254;
			7283: outdata = 32'd58253;
			7284: outdata = 32'd58252;
			7285: outdata = 32'd58251;
			7286: outdata = 32'd58250;
			7287: outdata = 32'd58249;
			7288: outdata = 32'd58248;
			7289: outdata = 32'd58247;
			7290: outdata = 32'd58246;
			7291: outdata = 32'd58245;
			7292: outdata = 32'd58244;
			7293: outdata = 32'd58243;
			7294: outdata = 32'd58242;
			7295: outdata = 32'd58241;
			7296: outdata = 32'd58240;
			7297: outdata = 32'd58239;
			7298: outdata = 32'd58238;
			7299: outdata = 32'd58237;
			7300: outdata = 32'd58236;
			7301: outdata = 32'd58235;
			7302: outdata = 32'd58234;
			7303: outdata = 32'd58233;
			7304: outdata = 32'd58232;
			7305: outdata = 32'd58231;
			7306: outdata = 32'd58230;
			7307: outdata = 32'd58229;
			7308: outdata = 32'd58228;
			7309: outdata = 32'd58227;
			7310: outdata = 32'd58226;
			7311: outdata = 32'd58225;
			7312: outdata = 32'd58224;
			7313: outdata = 32'd58223;
			7314: outdata = 32'd58222;
			7315: outdata = 32'd58221;
			7316: outdata = 32'd58220;
			7317: outdata = 32'd58219;
			7318: outdata = 32'd58218;
			7319: outdata = 32'd58217;
			7320: outdata = 32'd58216;
			7321: outdata = 32'd58215;
			7322: outdata = 32'd58214;
			7323: outdata = 32'd58213;
			7324: outdata = 32'd58212;
			7325: outdata = 32'd58211;
			7326: outdata = 32'd58210;
			7327: outdata = 32'd58209;
			7328: outdata = 32'd58208;
			7329: outdata = 32'd58207;
			7330: outdata = 32'd58206;
			7331: outdata = 32'd58205;
			7332: outdata = 32'd58204;
			7333: outdata = 32'd58203;
			7334: outdata = 32'd58202;
			7335: outdata = 32'd58201;
			7336: outdata = 32'd58200;
			7337: outdata = 32'd58199;
			7338: outdata = 32'd58198;
			7339: outdata = 32'd58197;
			7340: outdata = 32'd58196;
			7341: outdata = 32'd58195;
			7342: outdata = 32'd58194;
			7343: outdata = 32'd58193;
			7344: outdata = 32'd58192;
			7345: outdata = 32'd58191;
			7346: outdata = 32'd58190;
			7347: outdata = 32'd58189;
			7348: outdata = 32'd58188;
			7349: outdata = 32'd58187;
			7350: outdata = 32'd58186;
			7351: outdata = 32'd58185;
			7352: outdata = 32'd58184;
			7353: outdata = 32'd58183;
			7354: outdata = 32'd58182;
			7355: outdata = 32'd58181;
			7356: outdata = 32'd58180;
			7357: outdata = 32'd58179;
			7358: outdata = 32'd58178;
			7359: outdata = 32'd58177;
			7360: outdata = 32'd58176;
			7361: outdata = 32'd58175;
			7362: outdata = 32'd58174;
			7363: outdata = 32'd58173;
			7364: outdata = 32'd58172;
			7365: outdata = 32'd58171;
			7366: outdata = 32'd58170;
			7367: outdata = 32'd58169;
			7368: outdata = 32'd58168;
			7369: outdata = 32'd58167;
			7370: outdata = 32'd58166;
			7371: outdata = 32'd58165;
			7372: outdata = 32'd58164;
			7373: outdata = 32'd58163;
			7374: outdata = 32'd58162;
			7375: outdata = 32'd58161;
			7376: outdata = 32'd58160;
			7377: outdata = 32'd58159;
			7378: outdata = 32'd58158;
			7379: outdata = 32'd58157;
			7380: outdata = 32'd58156;
			7381: outdata = 32'd58155;
			7382: outdata = 32'd58154;
			7383: outdata = 32'd58153;
			7384: outdata = 32'd58152;
			7385: outdata = 32'd58151;
			7386: outdata = 32'd58150;
			7387: outdata = 32'd58149;
			7388: outdata = 32'd58148;
			7389: outdata = 32'd58147;
			7390: outdata = 32'd58146;
			7391: outdata = 32'd58145;
			7392: outdata = 32'd58144;
			7393: outdata = 32'd58143;
			7394: outdata = 32'd58142;
			7395: outdata = 32'd58141;
			7396: outdata = 32'd58140;
			7397: outdata = 32'd58139;
			7398: outdata = 32'd58138;
			7399: outdata = 32'd58137;
			7400: outdata = 32'd58136;
			7401: outdata = 32'd58135;
			7402: outdata = 32'd58134;
			7403: outdata = 32'd58133;
			7404: outdata = 32'd58132;
			7405: outdata = 32'd58131;
			7406: outdata = 32'd58130;
			7407: outdata = 32'd58129;
			7408: outdata = 32'd58128;
			7409: outdata = 32'd58127;
			7410: outdata = 32'd58126;
			7411: outdata = 32'd58125;
			7412: outdata = 32'd58124;
			7413: outdata = 32'd58123;
			7414: outdata = 32'd58122;
			7415: outdata = 32'd58121;
			7416: outdata = 32'd58120;
			7417: outdata = 32'd58119;
			7418: outdata = 32'd58118;
			7419: outdata = 32'd58117;
			7420: outdata = 32'd58116;
			7421: outdata = 32'd58115;
			7422: outdata = 32'd58114;
			7423: outdata = 32'd58113;
			7424: outdata = 32'd58112;
			7425: outdata = 32'd58111;
			7426: outdata = 32'd58110;
			7427: outdata = 32'd58109;
			7428: outdata = 32'd58108;
			7429: outdata = 32'd58107;
			7430: outdata = 32'd58106;
			7431: outdata = 32'd58105;
			7432: outdata = 32'd58104;
			7433: outdata = 32'd58103;
			7434: outdata = 32'd58102;
			7435: outdata = 32'd58101;
			7436: outdata = 32'd58100;
			7437: outdata = 32'd58099;
			7438: outdata = 32'd58098;
			7439: outdata = 32'd58097;
			7440: outdata = 32'd58096;
			7441: outdata = 32'd58095;
			7442: outdata = 32'd58094;
			7443: outdata = 32'd58093;
			7444: outdata = 32'd58092;
			7445: outdata = 32'd58091;
			7446: outdata = 32'd58090;
			7447: outdata = 32'd58089;
			7448: outdata = 32'd58088;
			7449: outdata = 32'd58087;
			7450: outdata = 32'd58086;
			7451: outdata = 32'd58085;
			7452: outdata = 32'd58084;
			7453: outdata = 32'd58083;
			7454: outdata = 32'd58082;
			7455: outdata = 32'd58081;
			7456: outdata = 32'd58080;
			7457: outdata = 32'd58079;
			7458: outdata = 32'd58078;
			7459: outdata = 32'd58077;
			7460: outdata = 32'd58076;
			7461: outdata = 32'd58075;
			7462: outdata = 32'd58074;
			7463: outdata = 32'd58073;
			7464: outdata = 32'd58072;
			7465: outdata = 32'd58071;
			7466: outdata = 32'd58070;
			7467: outdata = 32'd58069;
			7468: outdata = 32'd58068;
			7469: outdata = 32'd58067;
			7470: outdata = 32'd58066;
			7471: outdata = 32'd58065;
			7472: outdata = 32'd58064;
			7473: outdata = 32'd58063;
			7474: outdata = 32'd58062;
			7475: outdata = 32'd58061;
			7476: outdata = 32'd58060;
			7477: outdata = 32'd58059;
			7478: outdata = 32'd58058;
			7479: outdata = 32'd58057;
			7480: outdata = 32'd58056;
			7481: outdata = 32'd58055;
			7482: outdata = 32'd58054;
			7483: outdata = 32'd58053;
			7484: outdata = 32'd58052;
			7485: outdata = 32'd58051;
			7486: outdata = 32'd58050;
			7487: outdata = 32'd58049;
			7488: outdata = 32'd58048;
			7489: outdata = 32'd58047;
			7490: outdata = 32'd58046;
			7491: outdata = 32'd58045;
			7492: outdata = 32'd58044;
			7493: outdata = 32'd58043;
			7494: outdata = 32'd58042;
			7495: outdata = 32'd58041;
			7496: outdata = 32'd58040;
			7497: outdata = 32'd58039;
			7498: outdata = 32'd58038;
			7499: outdata = 32'd58037;
			7500: outdata = 32'd58036;
			7501: outdata = 32'd58035;
			7502: outdata = 32'd58034;
			7503: outdata = 32'd58033;
			7504: outdata = 32'd58032;
			7505: outdata = 32'd58031;
			7506: outdata = 32'd58030;
			7507: outdata = 32'd58029;
			7508: outdata = 32'd58028;
			7509: outdata = 32'd58027;
			7510: outdata = 32'd58026;
			7511: outdata = 32'd58025;
			7512: outdata = 32'd58024;
			7513: outdata = 32'd58023;
			7514: outdata = 32'd58022;
			7515: outdata = 32'd58021;
			7516: outdata = 32'd58020;
			7517: outdata = 32'd58019;
			7518: outdata = 32'd58018;
			7519: outdata = 32'd58017;
			7520: outdata = 32'd58016;
			7521: outdata = 32'd58015;
			7522: outdata = 32'd58014;
			7523: outdata = 32'd58013;
			7524: outdata = 32'd58012;
			7525: outdata = 32'd58011;
			7526: outdata = 32'd58010;
			7527: outdata = 32'd58009;
			7528: outdata = 32'd58008;
			7529: outdata = 32'd58007;
			7530: outdata = 32'd58006;
			7531: outdata = 32'd58005;
			7532: outdata = 32'd58004;
			7533: outdata = 32'd58003;
			7534: outdata = 32'd58002;
			7535: outdata = 32'd58001;
			7536: outdata = 32'd58000;
			7537: outdata = 32'd57999;
			7538: outdata = 32'd57998;
			7539: outdata = 32'd57997;
			7540: outdata = 32'd57996;
			7541: outdata = 32'd57995;
			7542: outdata = 32'd57994;
			7543: outdata = 32'd57993;
			7544: outdata = 32'd57992;
			7545: outdata = 32'd57991;
			7546: outdata = 32'd57990;
			7547: outdata = 32'd57989;
			7548: outdata = 32'd57988;
			7549: outdata = 32'd57987;
			7550: outdata = 32'd57986;
			7551: outdata = 32'd57985;
			7552: outdata = 32'd57984;
			7553: outdata = 32'd57983;
			7554: outdata = 32'd57982;
			7555: outdata = 32'd57981;
			7556: outdata = 32'd57980;
			7557: outdata = 32'd57979;
			7558: outdata = 32'd57978;
			7559: outdata = 32'd57977;
			7560: outdata = 32'd57976;
			7561: outdata = 32'd57975;
			7562: outdata = 32'd57974;
			7563: outdata = 32'd57973;
			7564: outdata = 32'd57972;
			7565: outdata = 32'd57971;
			7566: outdata = 32'd57970;
			7567: outdata = 32'd57969;
			7568: outdata = 32'd57968;
			7569: outdata = 32'd57967;
			7570: outdata = 32'd57966;
			7571: outdata = 32'd57965;
			7572: outdata = 32'd57964;
			7573: outdata = 32'd57963;
			7574: outdata = 32'd57962;
			7575: outdata = 32'd57961;
			7576: outdata = 32'd57960;
			7577: outdata = 32'd57959;
			7578: outdata = 32'd57958;
			7579: outdata = 32'd57957;
			7580: outdata = 32'd57956;
			7581: outdata = 32'd57955;
			7582: outdata = 32'd57954;
			7583: outdata = 32'd57953;
			7584: outdata = 32'd57952;
			7585: outdata = 32'd57951;
			7586: outdata = 32'd57950;
			7587: outdata = 32'd57949;
			7588: outdata = 32'd57948;
			7589: outdata = 32'd57947;
			7590: outdata = 32'd57946;
			7591: outdata = 32'd57945;
			7592: outdata = 32'd57944;
			7593: outdata = 32'd57943;
			7594: outdata = 32'd57942;
			7595: outdata = 32'd57941;
			7596: outdata = 32'd57940;
			7597: outdata = 32'd57939;
			7598: outdata = 32'd57938;
			7599: outdata = 32'd57937;
			7600: outdata = 32'd57936;
			7601: outdata = 32'd57935;
			7602: outdata = 32'd57934;
			7603: outdata = 32'd57933;
			7604: outdata = 32'd57932;
			7605: outdata = 32'd57931;
			7606: outdata = 32'd57930;
			7607: outdata = 32'd57929;
			7608: outdata = 32'd57928;
			7609: outdata = 32'd57927;
			7610: outdata = 32'd57926;
			7611: outdata = 32'd57925;
			7612: outdata = 32'd57924;
			7613: outdata = 32'd57923;
			7614: outdata = 32'd57922;
			7615: outdata = 32'd57921;
			7616: outdata = 32'd57920;
			7617: outdata = 32'd57919;
			7618: outdata = 32'd57918;
			7619: outdata = 32'd57917;
			7620: outdata = 32'd57916;
			7621: outdata = 32'd57915;
			7622: outdata = 32'd57914;
			7623: outdata = 32'd57913;
			7624: outdata = 32'd57912;
			7625: outdata = 32'd57911;
			7626: outdata = 32'd57910;
			7627: outdata = 32'd57909;
			7628: outdata = 32'd57908;
			7629: outdata = 32'd57907;
			7630: outdata = 32'd57906;
			7631: outdata = 32'd57905;
			7632: outdata = 32'd57904;
			7633: outdata = 32'd57903;
			7634: outdata = 32'd57902;
			7635: outdata = 32'd57901;
			7636: outdata = 32'd57900;
			7637: outdata = 32'd57899;
			7638: outdata = 32'd57898;
			7639: outdata = 32'd57897;
			7640: outdata = 32'd57896;
			7641: outdata = 32'd57895;
			7642: outdata = 32'd57894;
			7643: outdata = 32'd57893;
			7644: outdata = 32'd57892;
			7645: outdata = 32'd57891;
			7646: outdata = 32'd57890;
			7647: outdata = 32'd57889;
			7648: outdata = 32'd57888;
			7649: outdata = 32'd57887;
			7650: outdata = 32'd57886;
			7651: outdata = 32'd57885;
			7652: outdata = 32'd57884;
			7653: outdata = 32'd57883;
			7654: outdata = 32'd57882;
			7655: outdata = 32'd57881;
			7656: outdata = 32'd57880;
			7657: outdata = 32'd57879;
			7658: outdata = 32'd57878;
			7659: outdata = 32'd57877;
			7660: outdata = 32'd57876;
			7661: outdata = 32'd57875;
			7662: outdata = 32'd57874;
			7663: outdata = 32'd57873;
			7664: outdata = 32'd57872;
			7665: outdata = 32'd57871;
			7666: outdata = 32'd57870;
			7667: outdata = 32'd57869;
			7668: outdata = 32'd57868;
			7669: outdata = 32'd57867;
			7670: outdata = 32'd57866;
			7671: outdata = 32'd57865;
			7672: outdata = 32'd57864;
			7673: outdata = 32'd57863;
			7674: outdata = 32'd57862;
			7675: outdata = 32'd57861;
			7676: outdata = 32'd57860;
			7677: outdata = 32'd57859;
			7678: outdata = 32'd57858;
			7679: outdata = 32'd57857;
			7680: outdata = 32'd57856;
			7681: outdata = 32'd57855;
			7682: outdata = 32'd57854;
			7683: outdata = 32'd57853;
			7684: outdata = 32'd57852;
			7685: outdata = 32'd57851;
			7686: outdata = 32'd57850;
			7687: outdata = 32'd57849;
			7688: outdata = 32'd57848;
			7689: outdata = 32'd57847;
			7690: outdata = 32'd57846;
			7691: outdata = 32'd57845;
			7692: outdata = 32'd57844;
			7693: outdata = 32'd57843;
			7694: outdata = 32'd57842;
			7695: outdata = 32'd57841;
			7696: outdata = 32'd57840;
			7697: outdata = 32'd57839;
			7698: outdata = 32'd57838;
			7699: outdata = 32'd57837;
			7700: outdata = 32'd57836;
			7701: outdata = 32'd57835;
			7702: outdata = 32'd57834;
			7703: outdata = 32'd57833;
			7704: outdata = 32'd57832;
			7705: outdata = 32'd57831;
			7706: outdata = 32'd57830;
			7707: outdata = 32'd57829;
			7708: outdata = 32'd57828;
			7709: outdata = 32'd57827;
			7710: outdata = 32'd57826;
			7711: outdata = 32'd57825;
			7712: outdata = 32'd57824;
			7713: outdata = 32'd57823;
			7714: outdata = 32'd57822;
			7715: outdata = 32'd57821;
			7716: outdata = 32'd57820;
			7717: outdata = 32'd57819;
			7718: outdata = 32'd57818;
			7719: outdata = 32'd57817;
			7720: outdata = 32'd57816;
			7721: outdata = 32'd57815;
			7722: outdata = 32'd57814;
			7723: outdata = 32'd57813;
			7724: outdata = 32'd57812;
			7725: outdata = 32'd57811;
			7726: outdata = 32'd57810;
			7727: outdata = 32'd57809;
			7728: outdata = 32'd57808;
			7729: outdata = 32'd57807;
			7730: outdata = 32'd57806;
			7731: outdata = 32'd57805;
			7732: outdata = 32'd57804;
			7733: outdata = 32'd57803;
			7734: outdata = 32'd57802;
			7735: outdata = 32'd57801;
			7736: outdata = 32'd57800;
			7737: outdata = 32'd57799;
			7738: outdata = 32'd57798;
			7739: outdata = 32'd57797;
			7740: outdata = 32'd57796;
			7741: outdata = 32'd57795;
			7742: outdata = 32'd57794;
			7743: outdata = 32'd57793;
			7744: outdata = 32'd57792;
			7745: outdata = 32'd57791;
			7746: outdata = 32'd57790;
			7747: outdata = 32'd57789;
			7748: outdata = 32'd57788;
			7749: outdata = 32'd57787;
			7750: outdata = 32'd57786;
			7751: outdata = 32'd57785;
			7752: outdata = 32'd57784;
			7753: outdata = 32'd57783;
			7754: outdata = 32'd57782;
			7755: outdata = 32'd57781;
			7756: outdata = 32'd57780;
			7757: outdata = 32'd57779;
			7758: outdata = 32'd57778;
			7759: outdata = 32'd57777;
			7760: outdata = 32'd57776;
			7761: outdata = 32'd57775;
			7762: outdata = 32'd57774;
			7763: outdata = 32'd57773;
			7764: outdata = 32'd57772;
			7765: outdata = 32'd57771;
			7766: outdata = 32'd57770;
			7767: outdata = 32'd57769;
			7768: outdata = 32'd57768;
			7769: outdata = 32'd57767;
			7770: outdata = 32'd57766;
			7771: outdata = 32'd57765;
			7772: outdata = 32'd57764;
			7773: outdata = 32'd57763;
			7774: outdata = 32'd57762;
			7775: outdata = 32'd57761;
			7776: outdata = 32'd57760;
			7777: outdata = 32'd57759;
			7778: outdata = 32'd57758;
			7779: outdata = 32'd57757;
			7780: outdata = 32'd57756;
			7781: outdata = 32'd57755;
			7782: outdata = 32'd57754;
			7783: outdata = 32'd57753;
			7784: outdata = 32'd57752;
			7785: outdata = 32'd57751;
			7786: outdata = 32'd57750;
			7787: outdata = 32'd57749;
			7788: outdata = 32'd57748;
			7789: outdata = 32'd57747;
			7790: outdata = 32'd57746;
			7791: outdata = 32'd57745;
			7792: outdata = 32'd57744;
			7793: outdata = 32'd57743;
			7794: outdata = 32'd57742;
			7795: outdata = 32'd57741;
			7796: outdata = 32'd57740;
			7797: outdata = 32'd57739;
			7798: outdata = 32'd57738;
			7799: outdata = 32'd57737;
			7800: outdata = 32'd57736;
			7801: outdata = 32'd57735;
			7802: outdata = 32'd57734;
			7803: outdata = 32'd57733;
			7804: outdata = 32'd57732;
			7805: outdata = 32'd57731;
			7806: outdata = 32'd57730;
			7807: outdata = 32'd57729;
			7808: outdata = 32'd57728;
			7809: outdata = 32'd57727;
			7810: outdata = 32'd57726;
			7811: outdata = 32'd57725;
			7812: outdata = 32'd57724;
			7813: outdata = 32'd57723;
			7814: outdata = 32'd57722;
			7815: outdata = 32'd57721;
			7816: outdata = 32'd57720;
			7817: outdata = 32'd57719;
			7818: outdata = 32'd57718;
			7819: outdata = 32'd57717;
			7820: outdata = 32'd57716;
			7821: outdata = 32'd57715;
			7822: outdata = 32'd57714;
			7823: outdata = 32'd57713;
			7824: outdata = 32'd57712;
			7825: outdata = 32'd57711;
			7826: outdata = 32'd57710;
			7827: outdata = 32'd57709;
			7828: outdata = 32'd57708;
			7829: outdata = 32'd57707;
			7830: outdata = 32'd57706;
			7831: outdata = 32'd57705;
			7832: outdata = 32'd57704;
			7833: outdata = 32'd57703;
			7834: outdata = 32'd57702;
			7835: outdata = 32'd57701;
			7836: outdata = 32'd57700;
			7837: outdata = 32'd57699;
			7838: outdata = 32'd57698;
			7839: outdata = 32'd57697;
			7840: outdata = 32'd57696;
			7841: outdata = 32'd57695;
			7842: outdata = 32'd57694;
			7843: outdata = 32'd57693;
			7844: outdata = 32'd57692;
			7845: outdata = 32'd57691;
			7846: outdata = 32'd57690;
			7847: outdata = 32'd57689;
			7848: outdata = 32'd57688;
			7849: outdata = 32'd57687;
			7850: outdata = 32'd57686;
			7851: outdata = 32'd57685;
			7852: outdata = 32'd57684;
			7853: outdata = 32'd57683;
			7854: outdata = 32'd57682;
			7855: outdata = 32'd57681;
			7856: outdata = 32'd57680;
			7857: outdata = 32'd57679;
			7858: outdata = 32'd57678;
			7859: outdata = 32'd57677;
			7860: outdata = 32'd57676;
			7861: outdata = 32'd57675;
			7862: outdata = 32'd57674;
			7863: outdata = 32'd57673;
			7864: outdata = 32'd57672;
			7865: outdata = 32'd57671;
			7866: outdata = 32'd57670;
			7867: outdata = 32'd57669;
			7868: outdata = 32'd57668;
			7869: outdata = 32'd57667;
			7870: outdata = 32'd57666;
			7871: outdata = 32'd57665;
			7872: outdata = 32'd57664;
			7873: outdata = 32'd57663;
			7874: outdata = 32'd57662;
			7875: outdata = 32'd57661;
			7876: outdata = 32'd57660;
			7877: outdata = 32'd57659;
			7878: outdata = 32'd57658;
			7879: outdata = 32'd57657;
			7880: outdata = 32'd57656;
			7881: outdata = 32'd57655;
			7882: outdata = 32'd57654;
			7883: outdata = 32'd57653;
			7884: outdata = 32'd57652;
			7885: outdata = 32'd57651;
			7886: outdata = 32'd57650;
			7887: outdata = 32'd57649;
			7888: outdata = 32'd57648;
			7889: outdata = 32'd57647;
			7890: outdata = 32'd57646;
			7891: outdata = 32'd57645;
			7892: outdata = 32'd57644;
			7893: outdata = 32'd57643;
			7894: outdata = 32'd57642;
			7895: outdata = 32'd57641;
			7896: outdata = 32'd57640;
			7897: outdata = 32'd57639;
			7898: outdata = 32'd57638;
			7899: outdata = 32'd57637;
			7900: outdata = 32'd57636;
			7901: outdata = 32'd57635;
			7902: outdata = 32'd57634;
			7903: outdata = 32'd57633;
			7904: outdata = 32'd57632;
			7905: outdata = 32'd57631;
			7906: outdata = 32'd57630;
			7907: outdata = 32'd57629;
			7908: outdata = 32'd57628;
			7909: outdata = 32'd57627;
			7910: outdata = 32'd57626;
			7911: outdata = 32'd57625;
			7912: outdata = 32'd57624;
			7913: outdata = 32'd57623;
			7914: outdata = 32'd57622;
			7915: outdata = 32'd57621;
			7916: outdata = 32'd57620;
			7917: outdata = 32'd57619;
			7918: outdata = 32'd57618;
			7919: outdata = 32'd57617;
			7920: outdata = 32'd57616;
			7921: outdata = 32'd57615;
			7922: outdata = 32'd57614;
			7923: outdata = 32'd57613;
			7924: outdata = 32'd57612;
			7925: outdata = 32'd57611;
			7926: outdata = 32'd57610;
			7927: outdata = 32'd57609;
			7928: outdata = 32'd57608;
			7929: outdata = 32'd57607;
			7930: outdata = 32'd57606;
			7931: outdata = 32'd57605;
			7932: outdata = 32'd57604;
			7933: outdata = 32'd57603;
			7934: outdata = 32'd57602;
			7935: outdata = 32'd57601;
			7936: outdata = 32'd57600;
			7937: outdata = 32'd57599;
			7938: outdata = 32'd57598;
			7939: outdata = 32'd57597;
			7940: outdata = 32'd57596;
			7941: outdata = 32'd57595;
			7942: outdata = 32'd57594;
			7943: outdata = 32'd57593;
			7944: outdata = 32'd57592;
			7945: outdata = 32'd57591;
			7946: outdata = 32'd57590;
			7947: outdata = 32'd57589;
			7948: outdata = 32'd57588;
			7949: outdata = 32'd57587;
			7950: outdata = 32'd57586;
			7951: outdata = 32'd57585;
			7952: outdata = 32'd57584;
			7953: outdata = 32'd57583;
			7954: outdata = 32'd57582;
			7955: outdata = 32'd57581;
			7956: outdata = 32'd57580;
			7957: outdata = 32'd57579;
			7958: outdata = 32'd57578;
			7959: outdata = 32'd57577;
			7960: outdata = 32'd57576;
			7961: outdata = 32'd57575;
			7962: outdata = 32'd57574;
			7963: outdata = 32'd57573;
			7964: outdata = 32'd57572;
			7965: outdata = 32'd57571;
			7966: outdata = 32'd57570;
			7967: outdata = 32'd57569;
			7968: outdata = 32'd57568;
			7969: outdata = 32'd57567;
			7970: outdata = 32'd57566;
			7971: outdata = 32'd57565;
			7972: outdata = 32'd57564;
			7973: outdata = 32'd57563;
			7974: outdata = 32'd57562;
			7975: outdata = 32'd57561;
			7976: outdata = 32'd57560;
			7977: outdata = 32'd57559;
			7978: outdata = 32'd57558;
			7979: outdata = 32'd57557;
			7980: outdata = 32'd57556;
			7981: outdata = 32'd57555;
			7982: outdata = 32'd57554;
			7983: outdata = 32'd57553;
			7984: outdata = 32'd57552;
			7985: outdata = 32'd57551;
			7986: outdata = 32'd57550;
			7987: outdata = 32'd57549;
			7988: outdata = 32'd57548;
			7989: outdata = 32'd57547;
			7990: outdata = 32'd57546;
			7991: outdata = 32'd57545;
			7992: outdata = 32'd57544;
			7993: outdata = 32'd57543;
			7994: outdata = 32'd57542;
			7995: outdata = 32'd57541;
			7996: outdata = 32'd57540;
			7997: outdata = 32'd57539;
			7998: outdata = 32'd57538;
			7999: outdata = 32'd57537;
			8000: outdata = 32'd57536;
			8001: outdata = 32'd57535;
			8002: outdata = 32'd57534;
			8003: outdata = 32'd57533;
			8004: outdata = 32'd57532;
			8005: outdata = 32'd57531;
			8006: outdata = 32'd57530;
			8007: outdata = 32'd57529;
			8008: outdata = 32'd57528;
			8009: outdata = 32'd57527;
			8010: outdata = 32'd57526;
			8011: outdata = 32'd57525;
			8012: outdata = 32'd57524;
			8013: outdata = 32'd57523;
			8014: outdata = 32'd57522;
			8015: outdata = 32'd57521;
			8016: outdata = 32'd57520;
			8017: outdata = 32'd57519;
			8018: outdata = 32'd57518;
			8019: outdata = 32'd57517;
			8020: outdata = 32'd57516;
			8021: outdata = 32'd57515;
			8022: outdata = 32'd57514;
			8023: outdata = 32'd57513;
			8024: outdata = 32'd57512;
			8025: outdata = 32'd57511;
			8026: outdata = 32'd57510;
			8027: outdata = 32'd57509;
			8028: outdata = 32'd57508;
			8029: outdata = 32'd57507;
			8030: outdata = 32'd57506;
			8031: outdata = 32'd57505;
			8032: outdata = 32'd57504;
			8033: outdata = 32'd57503;
			8034: outdata = 32'd57502;
			8035: outdata = 32'd57501;
			8036: outdata = 32'd57500;
			8037: outdata = 32'd57499;
			8038: outdata = 32'd57498;
			8039: outdata = 32'd57497;
			8040: outdata = 32'd57496;
			8041: outdata = 32'd57495;
			8042: outdata = 32'd57494;
			8043: outdata = 32'd57493;
			8044: outdata = 32'd57492;
			8045: outdata = 32'd57491;
			8046: outdata = 32'd57490;
			8047: outdata = 32'd57489;
			8048: outdata = 32'd57488;
			8049: outdata = 32'd57487;
			8050: outdata = 32'd57486;
			8051: outdata = 32'd57485;
			8052: outdata = 32'd57484;
			8053: outdata = 32'd57483;
			8054: outdata = 32'd57482;
			8055: outdata = 32'd57481;
			8056: outdata = 32'd57480;
			8057: outdata = 32'd57479;
			8058: outdata = 32'd57478;
			8059: outdata = 32'd57477;
			8060: outdata = 32'd57476;
			8061: outdata = 32'd57475;
			8062: outdata = 32'd57474;
			8063: outdata = 32'd57473;
			8064: outdata = 32'd57472;
			8065: outdata = 32'd57471;
			8066: outdata = 32'd57470;
			8067: outdata = 32'd57469;
			8068: outdata = 32'd57468;
			8069: outdata = 32'd57467;
			8070: outdata = 32'd57466;
			8071: outdata = 32'd57465;
			8072: outdata = 32'd57464;
			8073: outdata = 32'd57463;
			8074: outdata = 32'd57462;
			8075: outdata = 32'd57461;
			8076: outdata = 32'd57460;
			8077: outdata = 32'd57459;
			8078: outdata = 32'd57458;
			8079: outdata = 32'd57457;
			8080: outdata = 32'd57456;
			8081: outdata = 32'd57455;
			8082: outdata = 32'd57454;
			8083: outdata = 32'd57453;
			8084: outdata = 32'd57452;
			8085: outdata = 32'd57451;
			8086: outdata = 32'd57450;
			8087: outdata = 32'd57449;
			8088: outdata = 32'd57448;
			8089: outdata = 32'd57447;
			8090: outdata = 32'd57446;
			8091: outdata = 32'd57445;
			8092: outdata = 32'd57444;
			8093: outdata = 32'd57443;
			8094: outdata = 32'd57442;
			8095: outdata = 32'd57441;
			8096: outdata = 32'd57440;
			8097: outdata = 32'd57439;
			8098: outdata = 32'd57438;
			8099: outdata = 32'd57437;
			8100: outdata = 32'd57436;
			8101: outdata = 32'd57435;
			8102: outdata = 32'd57434;
			8103: outdata = 32'd57433;
			8104: outdata = 32'd57432;
			8105: outdata = 32'd57431;
			8106: outdata = 32'd57430;
			8107: outdata = 32'd57429;
			8108: outdata = 32'd57428;
			8109: outdata = 32'd57427;
			8110: outdata = 32'd57426;
			8111: outdata = 32'd57425;
			8112: outdata = 32'd57424;
			8113: outdata = 32'd57423;
			8114: outdata = 32'd57422;
			8115: outdata = 32'd57421;
			8116: outdata = 32'd57420;
			8117: outdata = 32'd57419;
			8118: outdata = 32'd57418;
			8119: outdata = 32'd57417;
			8120: outdata = 32'd57416;
			8121: outdata = 32'd57415;
			8122: outdata = 32'd57414;
			8123: outdata = 32'd57413;
			8124: outdata = 32'd57412;
			8125: outdata = 32'd57411;
			8126: outdata = 32'd57410;
			8127: outdata = 32'd57409;
			8128: outdata = 32'd57408;
			8129: outdata = 32'd57407;
			8130: outdata = 32'd57406;
			8131: outdata = 32'd57405;
			8132: outdata = 32'd57404;
			8133: outdata = 32'd57403;
			8134: outdata = 32'd57402;
			8135: outdata = 32'd57401;
			8136: outdata = 32'd57400;
			8137: outdata = 32'd57399;
			8138: outdata = 32'd57398;
			8139: outdata = 32'd57397;
			8140: outdata = 32'd57396;
			8141: outdata = 32'd57395;
			8142: outdata = 32'd57394;
			8143: outdata = 32'd57393;
			8144: outdata = 32'd57392;
			8145: outdata = 32'd57391;
			8146: outdata = 32'd57390;
			8147: outdata = 32'd57389;
			8148: outdata = 32'd57388;
			8149: outdata = 32'd57387;
			8150: outdata = 32'd57386;
			8151: outdata = 32'd57385;
			8152: outdata = 32'd57384;
			8153: outdata = 32'd57383;
			8154: outdata = 32'd57382;
			8155: outdata = 32'd57381;
			8156: outdata = 32'd57380;
			8157: outdata = 32'd57379;
			8158: outdata = 32'd57378;
			8159: outdata = 32'd57377;
			8160: outdata = 32'd57376;
			8161: outdata = 32'd57375;
			8162: outdata = 32'd57374;
			8163: outdata = 32'd57373;
			8164: outdata = 32'd57372;
			8165: outdata = 32'd57371;
			8166: outdata = 32'd57370;
			8167: outdata = 32'd57369;
			8168: outdata = 32'd57368;
			8169: outdata = 32'd57367;
			8170: outdata = 32'd57366;
			8171: outdata = 32'd57365;
			8172: outdata = 32'd57364;
			8173: outdata = 32'd57363;
			8174: outdata = 32'd57362;
			8175: outdata = 32'd57361;
			8176: outdata = 32'd57360;
			8177: outdata = 32'd57359;
			8178: outdata = 32'd57358;
			8179: outdata = 32'd57357;
			8180: outdata = 32'd57356;
			8181: outdata = 32'd57355;
			8182: outdata = 32'd57354;
			8183: outdata = 32'd57353;
			8184: outdata = 32'd57352;
			8185: outdata = 32'd57351;
			8186: outdata = 32'd57350;
			8187: outdata = 32'd57349;
			8188: outdata = 32'd57348;
			8189: outdata = 32'd57347;
			8190: outdata = 32'd57346;
			8191: outdata = 32'd57345;
			8192: outdata = 32'd57344;
			8193: outdata = 32'd57343;
			8194: outdata = 32'd57342;
			8195: outdata = 32'd57341;
			8196: outdata = 32'd57340;
			8197: outdata = 32'd57339;
			8198: outdata = 32'd57338;
			8199: outdata = 32'd57337;
			8200: outdata = 32'd57336;
			8201: outdata = 32'd57335;
			8202: outdata = 32'd57334;
			8203: outdata = 32'd57333;
			8204: outdata = 32'd57332;
			8205: outdata = 32'd57331;
			8206: outdata = 32'd57330;
			8207: outdata = 32'd57329;
			8208: outdata = 32'd57328;
			8209: outdata = 32'd57327;
			8210: outdata = 32'd57326;
			8211: outdata = 32'd57325;
			8212: outdata = 32'd57324;
			8213: outdata = 32'd57323;
			8214: outdata = 32'd57322;
			8215: outdata = 32'd57321;
			8216: outdata = 32'd57320;
			8217: outdata = 32'd57319;
			8218: outdata = 32'd57318;
			8219: outdata = 32'd57317;
			8220: outdata = 32'd57316;
			8221: outdata = 32'd57315;
			8222: outdata = 32'd57314;
			8223: outdata = 32'd57313;
			8224: outdata = 32'd57312;
			8225: outdata = 32'd57311;
			8226: outdata = 32'd57310;
			8227: outdata = 32'd57309;
			8228: outdata = 32'd57308;
			8229: outdata = 32'd57307;
			8230: outdata = 32'd57306;
			8231: outdata = 32'd57305;
			8232: outdata = 32'd57304;
			8233: outdata = 32'd57303;
			8234: outdata = 32'd57302;
			8235: outdata = 32'd57301;
			8236: outdata = 32'd57300;
			8237: outdata = 32'd57299;
			8238: outdata = 32'd57298;
			8239: outdata = 32'd57297;
			8240: outdata = 32'd57296;
			8241: outdata = 32'd57295;
			8242: outdata = 32'd57294;
			8243: outdata = 32'd57293;
			8244: outdata = 32'd57292;
			8245: outdata = 32'd57291;
			8246: outdata = 32'd57290;
			8247: outdata = 32'd57289;
			8248: outdata = 32'd57288;
			8249: outdata = 32'd57287;
			8250: outdata = 32'd57286;
			8251: outdata = 32'd57285;
			8252: outdata = 32'd57284;
			8253: outdata = 32'd57283;
			8254: outdata = 32'd57282;
			8255: outdata = 32'd57281;
			8256: outdata = 32'd57280;
			8257: outdata = 32'd57279;
			8258: outdata = 32'd57278;
			8259: outdata = 32'd57277;
			8260: outdata = 32'd57276;
			8261: outdata = 32'd57275;
			8262: outdata = 32'd57274;
			8263: outdata = 32'd57273;
			8264: outdata = 32'd57272;
			8265: outdata = 32'd57271;
			8266: outdata = 32'd57270;
			8267: outdata = 32'd57269;
			8268: outdata = 32'd57268;
			8269: outdata = 32'd57267;
			8270: outdata = 32'd57266;
			8271: outdata = 32'd57265;
			8272: outdata = 32'd57264;
			8273: outdata = 32'd57263;
			8274: outdata = 32'd57262;
			8275: outdata = 32'd57261;
			8276: outdata = 32'd57260;
			8277: outdata = 32'd57259;
			8278: outdata = 32'd57258;
			8279: outdata = 32'd57257;
			8280: outdata = 32'd57256;
			8281: outdata = 32'd57255;
			8282: outdata = 32'd57254;
			8283: outdata = 32'd57253;
			8284: outdata = 32'd57252;
			8285: outdata = 32'd57251;
			8286: outdata = 32'd57250;
			8287: outdata = 32'd57249;
			8288: outdata = 32'd57248;
			8289: outdata = 32'd57247;
			8290: outdata = 32'd57246;
			8291: outdata = 32'd57245;
			8292: outdata = 32'd57244;
			8293: outdata = 32'd57243;
			8294: outdata = 32'd57242;
			8295: outdata = 32'd57241;
			8296: outdata = 32'd57240;
			8297: outdata = 32'd57239;
			8298: outdata = 32'd57238;
			8299: outdata = 32'd57237;
			8300: outdata = 32'd57236;
			8301: outdata = 32'd57235;
			8302: outdata = 32'd57234;
			8303: outdata = 32'd57233;
			8304: outdata = 32'd57232;
			8305: outdata = 32'd57231;
			8306: outdata = 32'd57230;
			8307: outdata = 32'd57229;
			8308: outdata = 32'd57228;
			8309: outdata = 32'd57227;
			8310: outdata = 32'd57226;
			8311: outdata = 32'd57225;
			8312: outdata = 32'd57224;
			8313: outdata = 32'd57223;
			8314: outdata = 32'd57222;
			8315: outdata = 32'd57221;
			8316: outdata = 32'd57220;
			8317: outdata = 32'd57219;
			8318: outdata = 32'd57218;
			8319: outdata = 32'd57217;
			8320: outdata = 32'd57216;
			8321: outdata = 32'd57215;
			8322: outdata = 32'd57214;
			8323: outdata = 32'd57213;
			8324: outdata = 32'd57212;
			8325: outdata = 32'd57211;
			8326: outdata = 32'd57210;
			8327: outdata = 32'd57209;
			8328: outdata = 32'd57208;
			8329: outdata = 32'd57207;
			8330: outdata = 32'd57206;
			8331: outdata = 32'd57205;
			8332: outdata = 32'd57204;
			8333: outdata = 32'd57203;
			8334: outdata = 32'd57202;
			8335: outdata = 32'd57201;
			8336: outdata = 32'd57200;
			8337: outdata = 32'd57199;
			8338: outdata = 32'd57198;
			8339: outdata = 32'd57197;
			8340: outdata = 32'd57196;
			8341: outdata = 32'd57195;
			8342: outdata = 32'd57194;
			8343: outdata = 32'd57193;
			8344: outdata = 32'd57192;
			8345: outdata = 32'd57191;
			8346: outdata = 32'd57190;
			8347: outdata = 32'd57189;
			8348: outdata = 32'd57188;
			8349: outdata = 32'd57187;
			8350: outdata = 32'd57186;
			8351: outdata = 32'd57185;
			8352: outdata = 32'd57184;
			8353: outdata = 32'd57183;
			8354: outdata = 32'd57182;
			8355: outdata = 32'd57181;
			8356: outdata = 32'd57180;
			8357: outdata = 32'd57179;
			8358: outdata = 32'd57178;
			8359: outdata = 32'd57177;
			8360: outdata = 32'd57176;
			8361: outdata = 32'd57175;
			8362: outdata = 32'd57174;
			8363: outdata = 32'd57173;
			8364: outdata = 32'd57172;
			8365: outdata = 32'd57171;
			8366: outdata = 32'd57170;
			8367: outdata = 32'd57169;
			8368: outdata = 32'd57168;
			8369: outdata = 32'd57167;
			8370: outdata = 32'd57166;
			8371: outdata = 32'd57165;
			8372: outdata = 32'd57164;
			8373: outdata = 32'd57163;
			8374: outdata = 32'd57162;
			8375: outdata = 32'd57161;
			8376: outdata = 32'd57160;
			8377: outdata = 32'd57159;
			8378: outdata = 32'd57158;
			8379: outdata = 32'd57157;
			8380: outdata = 32'd57156;
			8381: outdata = 32'd57155;
			8382: outdata = 32'd57154;
			8383: outdata = 32'd57153;
			8384: outdata = 32'd57152;
			8385: outdata = 32'd57151;
			8386: outdata = 32'd57150;
			8387: outdata = 32'd57149;
			8388: outdata = 32'd57148;
			8389: outdata = 32'd57147;
			8390: outdata = 32'd57146;
			8391: outdata = 32'd57145;
			8392: outdata = 32'd57144;
			8393: outdata = 32'd57143;
			8394: outdata = 32'd57142;
			8395: outdata = 32'd57141;
			8396: outdata = 32'd57140;
			8397: outdata = 32'd57139;
			8398: outdata = 32'd57138;
			8399: outdata = 32'd57137;
			8400: outdata = 32'd57136;
			8401: outdata = 32'd57135;
			8402: outdata = 32'd57134;
			8403: outdata = 32'd57133;
			8404: outdata = 32'd57132;
			8405: outdata = 32'd57131;
			8406: outdata = 32'd57130;
			8407: outdata = 32'd57129;
			8408: outdata = 32'd57128;
			8409: outdata = 32'd57127;
			8410: outdata = 32'd57126;
			8411: outdata = 32'd57125;
			8412: outdata = 32'd57124;
			8413: outdata = 32'd57123;
			8414: outdata = 32'd57122;
			8415: outdata = 32'd57121;
			8416: outdata = 32'd57120;
			8417: outdata = 32'd57119;
			8418: outdata = 32'd57118;
			8419: outdata = 32'd57117;
			8420: outdata = 32'd57116;
			8421: outdata = 32'd57115;
			8422: outdata = 32'd57114;
			8423: outdata = 32'd57113;
			8424: outdata = 32'd57112;
			8425: outdata = 32'd57111;
			8426: outdata = 32'd57110;
			8427: outdata = 32'd57109;
			8428: outdata = 32'd57108;
			8429: outdata = 32'd57107;
			8430: outdata = 32'd57106;
			8431: outdata = 32'd57105;
			8432: outdata = 32'd57104;
			8433: outdata = 32'd57103;
			8434: outdata = 32'd57102;
			8435: outdata = 32'd57101;
			8436: outdata = 32'd57100;
			8437: outdata = 32'd57099;
			8438: outdata = 32'd57098;
			8439: outdata = 32'd57097;
			8440: outdata = 32'd57096;
			8441: outdata = 32'd57095;
			8442: outdata = 32'd57094;
			8443: outdata = 32'd57093;
			8444: outdata = 32'd57092;
			8445: outdata = 32'd57091;
			8446: outdata = 32'd57090;
			8447: outdata = 32'd57089;
			8448: outdata = 32'd57088;
			8449: outdata = 32'd57087;
			8450: outdata = 32'd57086;
			8451: outdata = 32'd57085;
			8452: outdata = 32'd57084;
			8453: outdata = 32'd57083;
			8454: outdata = 32'd57082;
			8455: outdata = 32'd57081;
			8456: outdata = 32'd57080;
			8457: outdata = 32'd57079;
			8458: outdata = 32'd57078;
			8459: outdata = 32'd57077;
			8460: outdata = 32'd57076;
			8461: outdata = 32'd57075;
			8462: outdata = 32'd57074;
			8463: outdata = 32'd57073;
			8464: outdata = 32'd57072;
			8465: outdata = 32'd57071;
			8466: outdata = 32'd57070;
			8467: outdata = 32'd57069;
			8468: outdata = 32'd57068;
			8469: outdata = 32'd57067;
			8470: outdata = 32'd57066;
			8471: outdata = 32'd57065;
			8472: outdata = 32'd57064;
			8473: outdata = 32'd57063;
			8474: outdata = 32'd57062;
			8475: outdata = 32'd57061;
			8476: outdata = 32'd57060;
			8477: outdata = 32'd57059;
			8478: outdata = 32'd57058;
			8479: outdata = 32'd57057;
			8480: outdata = 32'd57056;
			8481: outdata = 32'd57055;
			8482: outdata = 32'd57054;
			8483: outdata = 32'd57053;
			8484: outdata = 32'd57052;
			8485: outdata = 32'd57051;
			8486: outdata = 32'd57050;
			8487: outdata = 32'd57049;
			8488: outdata = 32'd57048;
			8489: outdata = 32'd57047;
			8490: outdata = 32'd57046;
			8491: outdata = 32'd57045;
			8492: outdata = 32'd57044;
			8493: outdata = 32'd57043;
			8494: outdata = 32'd57042;
			8495: outdata = 32'd57041;
			8496: outdata = 32'd57040;
			8497: outdata = 32'd57039;
			8498: outdata = 32'd57038;
			8499: outdata = 32'd57037;
			8500: outdata = 32'd57036;
			8501: outdata = 32'd57035;
			8502: outdata = 32'd57034;
			8503: outdata = 32'd57033;
			8504: outdata = 32'd57032;
			8505: outdata = 32'd57031;
			8506: outdata = 32'd57030;
			8507: outdata = 32'd57029;
			8508: outdata = 32'd57028;
			8509: outdata = 32'd57027;
			8510: outdata = 32'd57026;
			8511: outdata = 32'd57025;
			8512: outdata = 32'd57024;
			8513: outdata = 32'd57023;
			8514: outdata = 32'd57022;
			8515: outdata = 32'd57021;
			8516: outdata = 32'd57020;
			8517: outdata = 32'd57019;
			8518: outdata = 32'd57018;
			8519: outdata = 32'd57017;
			8520: outdata = 32'd57016;
			8521: outdata = 32'd57015;
			8522: outdata = 32'd57014;
			8523: outdata = 32'd57013;
			8524: outdata = 32'd57012;
			8525: outdata = 32'd57011;
			8526: outdata = 32'd57010;
			8527: outdata = 32'd57009;
			8528: outdata = 32'd57008;
			8529: outdata = 32'd57007;
			8530: outdata = 32'd57006;
			8531: outdata = 32'd57005;
			8532: outdata = 32'd57004;
			8533: outdata = 32'd57003;
			8534: outdata = 32'd57002;
			8535: outdata = 32'd57001;
			8536: outdata = 32'd57000;
			8537: outdata = 32'd56999;
			8538: outdata = 32'd56998;
			8539: outdata = 32'd56997;
			8540: outdata = 32'd56996;
			8541: outdata = 32'd56995;
			8542: outdata = 32'd56994;
			8543: outdata = 32'd56993;
			8544: outdata = 32'd56992;
			8545: outdata = 32'd56991;
			8546: outdata = 32'd56990;
			8547: outdata = 32'd56989;
			8548: outdata = 32'd56988;
			8549: outdata = 32'd56987;
			8550: outdata = 32'd56986;
			8551: outdata = 32'd56985;
			8552: outdata = 32'd56984;
			8553: outdata = 32'd56983;
			8554: outdata = 32'd56982;
			8555: outdata = 32'd56981;
			8556: outdata = 32'd56980;
			8557: outdata = 32'd56979;
			8558: outdata = 32'd56978;
			8559: outdata = 32'd56977;
			8560: outdata = 32'd56976;
			8561: outdata = 32'd56975;
			8562: outdata = 32'd56974;
			8563: outdata = 32'd56973;
			8564: outdata = 32'd56972;
			8565: outdata = 32'd56971;
			8566: outdata = 32'd56970;
			8567: outdata = 32'd56969;
			8568: outdata = 32'd56968;
			8569: outdata = 32'd56967;
			8570: outdata = 32'd56966;
			8571: outdata = 32'd56965;
			8572: outdata = 32'd56964;
			8573: outdata = 32'd56963;
			8574: outdata = 32'd56962;
			8575: outdata = 32'd56961;
			8576: outdata = 32'd56960;
			8577: outdata = 32'd56959;
			8578: outdata = 32'd56958;
			8579: outdata = 32'd56957;
			8580: outdata = 32'd56956;
			8581: outdata = 32'd56955;
			8582: outdata = 32'd56954;
			8583: outdata = 32'd56953;
			8584: outdata = 32'd56952;
			8585: outdata = 32'd56951;
			8586: outdata = 32'd56950;
			8587: outdata = 32'd56949;
			8588: outdata = 32'd56948;
			8589: outdata = 32'd56947;
			8590: outdata = 32'd56946;
			8591: outdata = 32'd56945;
			8592: outdata = 32'd56944;
			8593: outdata = 32'd56943;
			8594: outdata = 32'd56942;
			8595: outdata = 32'd56941;
			8596: outdata = 32'd56940;
			8597: outdata = 32'd56939;
			8598: outdata = 32'd56938;
			8599: outdata = 32'd56937;
			8600: outdata = 32'd56936;
			8601: outdata = 32'd56935;
			8602: outdata = 32'd56934;
			8603: outdata = 32'd56933;
			8604: outdata = 32'd56932;
			8605: outdata = 32'd56931;
			8606: outdata = 32'd56930;
			8607: outdata = 32'd56929;
			8608: outdata = 32'd56928;
			8609: outdata = 32'd56927;
			8610: outdata = 32'd56926;
			8611: outdata = 32'd56925;
			8612: outdata = 32'd56924;
			8613: outdata = 32'd56923;
			8614: outdata = 32'd56922;
			8615: outdata = 32'd56921;
			8616: outdata = 32'd56920;
			8617: outdata = 32'd56919;
			8618: outdata = 32'd56918;
			8619: outdata = 32'd56917;
			8620: outdata = 32'd56916;
			8621: outdata = 32'd56915;
			8622: outdata = 32'd56914;
			8623: outdata = 32'd56913;
			8624: outdata = 32'd56912;
			8625: outdata = 32'd56911;
			8626: outdata = 32'd56910;
			8627: outdata = 32'd56909;
			8628: outdata = 32'd56908;
			8629: outdata = 32'd56907;
			8630: outdata = 32'd56906;
			8631: outdata = 32'd56905;
			8632: outdata = 32'd56904;
			8633: outdata = 32'd56903;
			8634: outdata = 32'd56902;
			8635: outdata = 32'd56901;
			8636: outdata = 32'd56900;
			8637: outdata = 32'd56899;
			8638: outdata = 32'd56898;
			8639: outdata = 32'd56897;
			8640: outdata = 32'd56896;
			8641: outdata = 32'd56895;
			8642: outdata = 32'd56894;
			8643: outdata = 32'd56893;
			8644: outdata = 32'd56892;
			8645: outdata = 32'd56891;
			8646: outdata = 32'd56890;
			8647: outdata = 32'd56889;
			8648: outdata = 32'd56888;
			8649: outdata = 32'd56887;
			8650: outdata = 32'd56886;
			8651: outdata = 32'd56885;
			8652: outdata = 32'd56884;
			8653: outdata = 32'd56883;
			8654: outdata = 32'd56882;
			8655: outdata = 32'd56881;
			8656: outdata = 32'd56880;
			8657: outdata = 32'd56879;
			8658: outdata = 32'd56878;
			8659: outdata = 32'd56877;
			8660: outdata = 32'd56876;
			8661: outdata = 32'd56875;
			8662: outdata = 32'd56874;
			8663: outdata = 32'd56873;
			8664: outdata = 32'd56872;
			8665: outdata = 32'd56871;
			8666: outdata = 32'd56870;
			8667: outdata = 32'd56869;
			8668: outdata = 32'd56868;
			8669: outdata = 32'd56867;
			8670: outdata = 32'd56866;
			8671: outdata = 32'd56865;
			8672: outdata = 32'd56864;
			8673: outdata = 32'd56863;
			8674: outdata = 32'd56862;
			8675: outdata = 32'd56861;
			8676: outdata = 32'd56860;
			8677: outdata = 32'd56859;
			8678: outdata = 32'd56858;
			8679: outdata = 32'd56857;
			8680: outdata = 32'd56856;
			8681: outdata = 32'd56855;
			8682: outdata = 32'd56854;
			8683: outdata = 32'd56853;
			8684: outdata = 32'd56852;
			8685: outdata = 32'd56851;
			8686: outdata = 32'd56850;
			8687: outdata = 32'd56849;
			8688: outdata = 32'd56848;
			8689: outdata = 32'd56847;
			8690: outdata = 32'd56846;
			8691: outdata = 32'd56845;
			8692: outdata = 32'd56844;
			8693: outdata = 32'd56843;
			8694: outdata = 32'd56842;
			8695: outdata = 32'd56841;
			8696: outdata = 32'd56840;
			8697: outdata = 32'd56839;
			8698: outdata = 32'd56838;
			8699: outdata = 32'd56837;
			8700: outdata = 32'd56836;
			8701: outdata = 32'd56835;
			8702: outdata = 32'd56834;
			8703: outdata = 32'd56833;
			8704: outdata = 32'd56832;
			8705: outdata = 32'd56831;
			8706: outdata = 32'd56830;
			8707: outdata = 32'd56829;
			8708: outdata = 32'd56828;
			8709: outdata = 32'd56827;
			8710: outdata = 32'd56826;
			8711: outdata = 32'd56825;
			8712: outdata = 32'd56824;
			8713: outdata = 32'd56823;
			8714: outdata = 32'd56822;
			8715: outdata = 32'd56821;
			8716: outdata = 32'd56820;
			8717: outdata = 32'd56819;
			8718: outdata = 32'd56818;
			8719: outdata = 32'd56817;
			8720: outdata = 32'd56816;
			8721: outdata = 32'd56815;
			8722: outdata = 32'd56814;
			8723: outdata = 32'd56813;
			8724: outdata = 32'd56812;
			8725: outdata = 32'd56811;
			8726: outdata = 32'd56810;
			8727: outdata = 32'd56809;
			8728: outdata = 32'd56808;
			8729: outdata = 32'd56807;
			8730: outdata = 32'd56806;
			8731: outdata = 32'd56805;
			8732: outdata = 32'd56804;
			8733: outdata = 32'd56803;
			8734: outdata = 32'd56802;
			8735: outdata = 32'd56801;
			8736: outdata = 32'd56800;
			8737: outdata = 32'd56799;
			8738: outdata = 32'd56798;
			8739: outdata = 32'd56797;
			8740: outdata = 32'd56796;
			8741: outdata = 32'd56795;
			8742: outdata = 32'd56794;
			8743: outdata = 32'd56793;
			8744: outdata = 32'd56792;
			8745: outdata = 32'd56791;
			8746: outdata = 32'd56790;
			8747: outdata = 32'd56789;
			8748: outdata = 32'd56788;
			8749: outdata = 32'd56787;
			8750: outdata = 32'd56786;
			8751: outdata = 32'd56785;
			8752: outdata = 32'd56784;
			8753: outdata = 32'd56783;
			8754: outdata = 32'd56782;
			8755: outdata = 32'd56781;
			8756: outdata = 32'd56780;
			8757: outdata = 32'd56779;
			8758: outdata = 32'd56778;
			8759: outdata = 32'd56777;
			8760: outdata = 32'd56776;
			8761: outdata = 32'd56775;
			8762: outdata = 32'd56774;
			8763: outdata = 32'd56773;
			8764: outdata = 32'd56772;
			8765: outdata = 32'd56771;
			8766: outdata = 32'd56770;
			8767: outdata = 32'd56769;
			8768: outdata = 32'd56768;
			8769: outdata = 32'd56767;
			8770: outdata = 32'd56766;
			8771: outdata = 32'd56765;
			8772: outdata = 32'd56764;
			8773: outdata = 32'd56763;
			8774: outdata = 32'd56762;
			8775: outdata = 32'd56761;
			8776: outdata = 32'd56760;
			8777: outdata = 32'd56759;
			8778: outdata = 32'd56758;
			8779: outdata = 32'd56757;
			8780: outdata = 32'd56756;
			8781: outdata = 32'd56755;
			8782: outdata = 32'd56754;
			8783: outdata = 32'd56753;
			8784: outdata = 32'd56752;
			8785: outdata = 32'd56751;
			8786: outdata = 32'd56750;
			8787: outdata = 32'd56749;
			8788: outdata = 32'd56748;
			8789: outdata = 32'd56747;
			8790: outdata = 32'd56746;
			8791: outdata = 32'd56745;
			8792: outdata = 32'd56744;
			8793: outdata = 32'd56743;
			8794: outdata = 32'd56742;
			8795: outdata = 32'd56741;
			8796: outdata = 32'd56740;
			8797: outdata = 32'd56739;
			8798: outdata = 32'd56738;
			8799: outdata = 32'd56737;
			8800: outdata = 32'd56736;
			8801: outdata = 32'd56735;
			8802: outdata = 32'd56734;
			8803: outdata = 32'd56733;
			8804: outdata = 32'd56732;
			8805: outdata = 32'd56731;
			8806: outdata = 32'd56730;
			8807: outdata = 32'd56729;
			8808: outdata = 32'd56728;
			8809: outdata = 32'd56727;
			8810: outdata = 32'd56726;
			8811: outdata = 32'd56725;
			8812: outdata = 32'd56724;
			8813: outdata = 32'd56723;
			8814: outdata = 32'd56722;
			8815: outdata = 32'd56721;
			8816: outdata = 32'd56720;
			8817: outdata = 32'd56719;
			8818: outdata = 32'd56718;
			8819: outdata = 32'd56717;
			8820: outdata = 32'd56716;
			8821: outdata = 32'd56715;
			8822: outdata = 32'd56714;
			8823: outdata = 32'd56713;
			8824: outdata = 32'd56712;
			8825: outdata = 32'd56711;
			8826: outdata = 32'd56710;
			8827: outdata = 32'd56709;
			8828: outdata = 32'd56708;
			8829: outdata = 32'd56707;
			8830: outdata = 32'd56706;
			8831: outdata = 32'd56705;
			8832: outdata = 32'd56704;
			8833: outdata = 32'd56703;
			8834: outdata = 32'd56702;
			8835: outdata = 32'd56701;
			8836: outdata = 32'd56700;
			8837: outdata = 32'd56699;
			8838: outdata = 32'd56698;
			8839: outdata = 32'd56697;
			8840: outdata = 32'd56696;
			8841: outdata = 32'd56695;
			8842: outdata = 32'd56694;
			8843: outdata = 32'd56693;
			8844: outdata = 32'd56692;
			8845: outdata = 32'd56691;
			8846: outdata = 32'd56690;
			8847: outdata = 32'd56689;
			8848: outdata = 32'd56688;
			8849: outdata = 32'd56687;
			8850: outdata = 32'd56686;
			8851: outdata = 32'd56685;
			8852: outdata = 32'd56684;
			8853: outdata = 32'd56683;
			8854: outdata = 32'd56682;
			8855: outdata = 32'd56681;
			8856: outdata = 32'd56680;
			8857: outdata = 32'd56679;
			8858: outdata = 32'd56678;
			8859: outdata = 32'd56677;
			8860: outdata = 32'd56676;
			8861: outdata = 32'd56675;
			8862: outdata = 32'd56674;
			8863: outdata = 32'd56673;
			8864: outdata = 32'd56672;
			8865: outdata = 32'd56671;
			8866: outdata = 32'd56670;
			8867: outdata = 32'd56669;
			8868: outdata = 32'd56668;
			8869: outdata = 32'd56667;
			8870: outdata = 32'd56666;
			8871: outdata = 32'd56665;
			8872: outdata = 32'd56664;
			8873: outdata = 32'd56663;
			8874: outdata = 32'd56662;
			8875: outdata = 32'd56661;
			8876: outdata = 32'd56660;
			8877: outdata = 32'd56659;
			8878: outdata = 32'd56658;
			8879: outdata = 32'd56657;
			8880: outdata = 32'd56656;
			8881: outdata = 32'd56655;
			8882: outdata = 32'd56654;
			8883: outdata = 32'd56653;
			8884: outdata = 32'd56652;
			8885: outdata = 32'd56651;
			8886: outdata = 32'd56650;
			8887: outdata = 32'd56649;
			8888: outdata = 32'd56648;
			8889: outdata = 32'd56647;
			8890: outdata = 32'd56646;
			8891: outdata = 32'd56645;
			8892: outdata = 32'd56644;
			8893: outdata = 32'd56643;
			8894: outdata = 32'd56642;
			8895: outdata = 32'd56641;
			8896: outdata = 32'd56640;
			8897: outdata = 32'd56639;
			8898: outdata = 32'd56638;
			8899: outdata = 32'd56637;
			8900: outdata = 32'd56636;
			8901: outdata = 32'd56635;
			8902: outdata = 32'd56634;
			8903: outdata = 32'd56633;
			8904: outdata = 32'd56632;
			8905: outdata = 32'd56631;
			8906: outdata = 32'd56630;
			8907: outdata = 32'd56629;
			8908: outdata = 32'd56628;
			8909: outdata = 32'd56627;
			8910: outdata = 32'd56626;
			8911: outdata = 32'd56625;
			8912: outdata = 32'd56624;
			8913: outdata = 32'd56623;
			8914: outdata = 32'd56622;
			8915: outdata = 32'd56621;
			8916: outdata = 32'd56620;
			8917: outdata = 32'd56619;
			8918: outdata = 32'd56618;
			8919: outdata = 32'd56617;
			8920: outdata = 32'd56616;
			8921: outdata = 32'd56615;
			8922: outdata = 32'd56614;
			8923: outdata = 32'd56613;
			8924: outdata = 32'd56612;
			8925: outdata = 32'd56611;
			8926: outdata = 32'd56610;
			8927: outdata = 32'd56609;
			8928: outdata = 32'd56608;
			8929: outdata = 32'd56607;
			8930: outdata = 32'd56606;
			8931: outdata = 32'd56605;
			8932: outdata = 32'd56604;
			8933: outdata = 32'd56603;
			8934: outdata = 32'd56602;
			8935: outdata = 32'd56601;
			8936: outdata = 32'd56600;
			8937: outdata = 32'd56599;
			8938: outdata = 32'd56598;
			8939: outdata = 32'd56597;
			8940: outdata = 32'd56596;
			8941: outdata = 32'd56595;
			8942: outdata = 32'd56594;
			8943: outdata = 32'd56593;
			8944: outdata = 32'd56592;
			8945: outdata = 32'd56591;
			8946: outdata = 32'd56590;
			8947: outdata = 32'd56589;
			8948: outdata = 32'd56588;
			8949: outdata = 32'd56587;
			8950: outdata = 32'd56586;
			8951: outdata = 32'd56585;
			8952: outdata = 32'd56584;
			8953: outdata = 32'd56583;
			8954: outdata = 32'd56582;
			8955: outdata = 32'd56581;
			8956: outdata = 32'd56580;
			8957: outdata = 32'd56579;
			8958: outdata = 32'd56578;
			8959: outdata = 32'd56577;
			8960: outdata = 32'd56576;
			8961: outdata = 32'd56575;
			8962: outdata = 32'd56574;
			8963: outdata = 32'd56573;
			8964: outdata = 32'd56572;
			8965: outdata = 32'd56571;
			8966: outdata = 32'd56570;
			8967: outdata = 32'd56569;
			8968: outdata = 32'd56568;
			8969: outdata = 32'd56567;
			8970: outdata = 32'd56566;
			8971: outdata = 32'd56565;
			8972: outdata = 32'd56564;
			8973: outdata = 32'd56563;
			8974: outdata = 32'd56562;
			8975: outdata = 32'd56561;
			8976: outdata = 32'd56560;
			8977: outdata = 32'd56559;
			8978: outdata = 32'd56558;
			8979: outdata = 32'd56557;
			8980: outdata = 32'd56556;
			8981: outdata = 32'd56555;
			8982: outdata = 32'd56554;
			8983: outdata = 32'd56553;
			8984: outdata = 32'd56552;
			8985: outdata = 32'd56551;
			8986: outdata = 32'd56550;
			8987: outdata = 32'd56549;
			8988: outdata = 32'd56548;
			8989: outdata = 32'd56547;
			8990: outdata = 32'd56546;
			8991: outdata = 32'd56545;
			8992: outdata = 32'd56544;
			8993: outdata = 32'd56543;
			8994: outdata = 32'd56542;
			8995: outdata = 32'd56541;
			8996: outdata = 32'd56540;
			8997: outdata = 32'd56539;
			8998: outdata = 32'd56538;
			8999: outdata = 32'd56537;
			9000: outdata = 32'd56536;
			9001: outdata = 32'd56535;
			9002: outdata = 32'd56534;
			9003: outdata = 32'd56533;
			9004: outdata = 32'd56532;
			9005: outdata = 32'd56531;
			9006: outdata = 32'd56530;
			9007: outdata = 32'd56529;
			9008: outdata = 32'd56528;
			9009: outdata = 32'd56527;
			9010: outdata = 32'd56526;
			9011: outdata = 32'd56525;
			9012: outdata = 32'd56524;
			9013: outdata = 32'd56523;
			9014: outdata = 32'd56522;
			9015: outdata = 32'd56521;
			9016: outdata = 32'd56520;
			9017: outdata = 32'd56519;
			9018: outdata = 32'd56518;
			9019: outdata = 32'd56517;
			9020: outdata = 32'd56516;
			9021: outdata = 32'd56515;
			9022: outdata = 32'd56514;
			9023: outdata = 32'd56513;
			9024: outdata = 32'd56512;
			9025: outdata = 32'd56511;
			9026: outdata = 32'd56510;
			9027: outdata = 32'd56509;
			9028: outdata = 32'd56508;
			9029: outdata = 32'd56507;
			9030: outdata = 32'd56506;
			9031: outdata = 32'd56505;
			9032: outdata = 32'd56504;
			9033: outdata = 32'd56503;
			9034: outdata = 32'd56502;
			9035: outdata = 32'd56501;
			9036: outdata = 32'd56500;
			9037: outdata = 32'd56499;
			9038: outdata = 32'd56498;
			9039: outdata = 32'd56497;
			9040: outdata = 32'd56496;
			9041: outdata = 32'd56495;
			9042: outdata = 32'd56494;
			9043: outdata = 32'd56493;
			9044: outdata = 32'd56492;
			9045: outdata = 32'd56491;
			9046: outdata = 32'd56490;
			9047: outdata = 32'd56489;
			9048: outdata = 32'd56488;
			9049: outdata = 32'd56487;
			9050: outdata = 32'd56486;
			9051: outdata = 32'd56485;
			9052: outdata = 32'd56484;
			9053: outdata = 32'd56483;
			9054: outdata = 32'd56482;
			9055: outdata = 32'd56481;
			9056: outdata = 32'd56480;
			9057: outdata = 32'd56479;
			9058: outdata = 32'd56478;
			9059: outdata = 32'd56477;
			9060: outdata = 32'd56476;
			9061: outdata = 32'd56475;
			9062: outdata = 32'd56474;
			9063: outdata = 32'd56473;
			9064: outdata = 32'd56472;
			9065: outdata = 32'd56471;
			9066: outdata = 32'd56470;
			9067: outdata = 32'd56469;
			9068: outdata = 32'd56468;
			9069: outdata = 32'd56467;
			9070: outdata = 32'd56466;
			9071: outdata = 32'd56465;
			9072: outdata = 32'd56464;
			9073: outdata = 32'd56463;
			9074: outdata = 32'd56462;
			9075: outdata = 32'd56461;
			9076: outdata = 32'd56460;
			9077: outdata = 32'd56459;
			9078: outdata = 32'd56458;
			9079: outdata = 32'd56457;
			9080: outdata = 32'd56456;
			9081: outdata = 32'd56455;
			9082: outdata = 32'd56454;
			9083: outdata = 32'd56453;
			9084: outdata = 32'd56452;
			9085: outdata = 32'd56451;
			9086: outdata = 32'd56450;
			9087: outdata = 32'd56449;
			9088: outdata = 32'd56448;
			9089: outdata = 32'd56447;
			9090: outdata = 32'd56446;
			9091: outdata = 32'd56445;
			9092: outdata = 32'd56444;
			9093: outdata = 32'd56443;
			9094: outdata = 32'd56442;
			9095: outdata = 32'd56441;
			9096: outdata = 32'd56440;
			9097: outdata = 32'd56439;
			9098: outdata = 32'd56438;
			9099: outdata = 32'd56437;
			9100: outdata = 32'd56436;
			9101: outdata = 32'd56435;
			9102: outdata = 32'd56434;
			9103: outdata = 32'd56433;
			9104: outdata = 32'd56432;
			9105: outdata = 32'd56431;
			9106: outdata = 32'd56430;
			9107: outdata = 32'd56429;
			9108: outdata = 32'd56428;
			9109: outdata = 32'd56427;
			9110: outdata = 32'd56426;
			9111: outdata = 32'd56425;
			9112: outdata = 32'd56424;
			9113: outdata = 32'd56423;
			9114: outdata = 32'd56422;
			9115: outdata = 32'd56421;
			9116: outdata = 32'd56420;
			9117: outdata = 32'd56419;
			9118: outdata = 32'd56418;
			9119: outdata = 32'd56417;
			9120: outdata = 32'd56416;
			9121: outdata = 32'd56415;
			9122: outdata = 32'd56414;
			9123: outdata = 32'd56413;
			9124: outdata = 32'd56412;
			9125: outdata = 32'd56411;
			9126: outdata = 32'd56410;
			9127: outdata = 32'd56409;
			9128: outdata = 32'd56408;
			9129: outdata = 32'd56407;
			9130: outdata = 32'd56406;
			9131: outdata = 32'd56405;
			9132: outdata = 32'd56404;
			9133: outdata = 32'd56403;
			9134: outdata = 32'd56402;
			9135: outdata = 32'd56401;
			9136: outdata = 32'd56400;
			9137: outdata = 32'd56399;
			9138: outdata = 32'd56398;
			9139: outdata = 32'd56397;
			9140: outdata = 32'd56396;
			9141: outdata = 32'd56395;
			9142: outdata = 32'd56394;
			9143: outdata = 32'd56393;
			9144: outdata = 32'd56392;
			9145: outdata = 32'd56391;
			9146: outdata = 32'd56390;
			9147: outdata = 32'd56389;
			9148: outdata = 32'd56388;
			9149: outdata = 32'd56387;
			9150: outdata = 32'd56386;
			9151: outdata = 32'd56385;
			9152: outdata = 32'd56384;
			9153: outdata = 32'd56383;
			9154: outdata = 32'd56382;
			9155: outdata = 32'd56381;
			9156: outdata = 32'd56380;
			9157: outdata = 32'd56379;
			9158: outdata = 32'd56378;
			9159: outdata = 32'd56377;
			9160: outdata = 32'd56376;
			9161: outdata = 32'd56375;
			9162: outdata = 32'd56374;
			9163: outdata = 32'd56373;
			9164: outdata = 32'd56372;
			9165: outdata = 32'd56371;
			9166: outdata = 32'd56370;
			9167: outdata = 32'd56369;
			9168: outdata = 32'd56368;
			9169: outdata = 32'd56367;
			9170: outdata = 32'd56366;
			9171: outdata = 32'd56365;
			9172: outdata = 32'd56364;
			9173: outdata = 32'd56363;
			9174: outdata = 32'd56362;
			9175: outdata = 32'd56361;
			9176: outdata = 32'd56360;
			9177: outdata = 32'd56359;
			9178: outdata = 32'd56358;
			9179: outdata = 32'd56357;
			9180: outdata = 32'd56356;
			9181: outdata = 32'd56355;
			9182: outdata = 32'd56354;
			9183: outdata = 32'd56353;
			9184: outdata = 32'd56352;
			9185: outdata = 32'd56351;
			9186: outdata = 32'd56350;
			9187: outdata = 32'd56349;
			9188: outdata = 32'd56348;
			9189: outdata = 32'd56347;
			9190: outdata = 32'd56346;
			9191: outdata = 32'd56345;
			9192: outdata = 32'd56344;
			9193: outdata = 32'd56343;
			9194: outdata = 32'd56342;
			9195: outdata = 32'd56341;
			9196: outdata = 32'd56340;
			9197: outdata = 32'd56339;
			9198: outdata = 32'd56338;
			9199: outdata = 32'd56337;
			9200: outdata = 32'd56336;
			9201: outdata = 32'd56335;
			9202: outdata = 32'd56334;
			9203: outdata = 32'd56333;
			9204: outdata = 32'd56332;
			9205: outdata = 32'd56331;
			9206: outdata = 32'd56330;
			9207: outdata = 32'd56329;
			9208: outdata = 32'd56328;
			9209: outdata = 32'd56327;
			9210: outdata = 32'd56326;
			9211: outdata = 32'd56325;
			9212: outdata = 32'd56324;
			9213: outdata = 32'd56323;
			9214: outdata = 32'd56322;
			9215: outdata = 32'd56321;
			9216: outdata = 32'd56320;
			9217: outdata = 32'd56319;
			9218: outdata = 32'd56318;
			9219: outdata = 32'd56317;
			9220: outdata = 32'd56316;
			9221: outdata = 32'd56315;
			9222: outdata = 32'd56314;
			9223: outdata = 32'd56313;
			9224: outdata = 32'd56312;
			9225: outdata = 32'd56311;
			9226: outdata = 32'd56310;
			9227: outdata = 32'd56309;
			9228: outdata = 32'd56308;
			9229: outdata = 32'd56307;
			9230: outdata = 32'd56306;
			9231: outdata = 32'd56305;
			9232: outdata = 32'd56304;
			9233: outdata = 32'd56303;
			9234: outdata = 32'd56302;
			9235: outdata = 32'd56301;
			9236: outdata = 32'd56300;
			9237: outdata = 32'd56299;
			9238: outdata = 32'd56298;
			9239: outdata = 32'd56297;
			9240: outdata = 32'd56296;
			9241: outdata = 32'd56295;
			9242: outdata = 32'd56294;
			9243: outdata = 32'd56293;
			9244: outdata = 32'd56292;
			9245: outdata = 32'd56291;
			9246: outdata = 32'd56290;
			9247: outdata = 32'd56289;
			9248: outdata = 32'd56288;
			9249: outdata = 32'd56287;
			9250: outdata = 32'd56286;
			9251: outdata = 32'd56285;
			9252: outdata = 32'd56284;
			9253: outdata = 32'd56283;
			9254: outdata = 32'd56282;
			9255: outdata = 32'd56281;
			9256: outdata = 32'd56280;
			9257: outdata = 32'd56279;
			9258: outdata = 32'd56278;
			9259: outdata = 32'd56277;
			9260: outdata = 32'd56276;
			9261: outdata = 32'd56275;
			9262: outdata = 32'd56274;
			9263: outdata = 32'd56273;
			9264: outdata = 32'd56272;
			9265: outdata = 32'd56271;
			9266: outdata = 32'd56270;
			9267: outdata = 32'd56269;
			9268: outdata = 32'd56268;
			9269: outdata = 32'd56267;
			9270: outdata = 32'd56266;
			9271: outdata = 32'd56265;
			9272: outdata = 32'd56264;
			9273: outdata = 32'd56263;
			9274: outdata = 32'd56262;
			9275: outdata = 32'd56261;
			9276: outdata = 32'd56260;
			9277: outdata = 32'd56259;
			9278: outdata = 32'd56258;
			9279: outdata = 32'd56257;
			9280: outdata = 32'd56256;
			9281: outdata = 32'd56255;
			9282: outdata = 32'd56254;
			9283: outdata = 32'd56253;
			9284: outdata = 32'd56252;
			9285: outdata = 32'd56251;
			9286: outdata = 32'd56250;
			9287: outdata = 32'd56249;
			9288: outdata = 32'd56248;
			9289: outdata = 32'd56247;
			9290: outdata = 32'd56246;
			9291: outdata = 32'd56245;
			9292: outdata = 32'd56244;
			9293: outdata = 32'd56243;
			9294: outdata = 32'd56242;
			9295: outdata = 32'd56241;
			9296: outdata = 32'd56240;
			9297: outdata = 32'd56239;
			9298: outdata = 32'd56238;
			9299: outdata = 32'd56237;
			9300: outdata = 32'd56236;
			9301: outdata = 32'd56235;
			9302: outdata = 32'd56234;
			9303: outdata = 32'd56233;
			9304: outdata = 32'd56232;
			9305: outdata = 32'd56231;
			9306: outdata = 32'd56230;
			9307: outdata = 32'd56229;
			9308: outdata = 32'd56228;
			9309: outdata = 32'd56227;
			9310: outdata = 32'd56226;
			9311: outdata = 32'd56225;
			9312: outdata = 32'd56224;
			9313: outdata = 32'd56223;
			9314: outdata = 32'd56222;
			9315: outdata = 32'd56221;
			9316: outdata = 32'd56220;
			9317: outdata = 32'd56219;
			9318: outdata = 32'd56218;
			9319: outdata = 32'd56217;
			9320: outdata = 32'd56216;
			9321: outdata = 32'd56215;
			9322: outdata = 32'd56214;
			9323: outdata = 32'd56213;
			9324: outdata = 32'd56212;
			9325: outdata = 32'd56211;
			9326: outdata = 32'd56210;
			9327: outdata = 32'd56209;
			9328: outdata = 32'd56208;
			9329: outdata = 32'd56207;
			9330: outdata = 32'd56206;
			9331: outdata = 32'd56205;
			9332: outdata = 32'd56204;
			9333: outdata = 32'd56203;
			9334: outdata = 32'd56202;
			9335: outdata = 32'd56201;
			9336: outdata = 32'd56200;
			9337: outdata = 32'd56199;
			9338: outdata = 32'd56198;
			9339: outdata = 32'd56197;
			9340: outdata = 32'd56196;
			9341: outdata = 32'd56195;
			9342: outdata = 32'd56194;
			9343: outdata = 32'd56193;
			9344: outdata = 32'd56192;
			9345: outdata = 32'd56191;
			9346: outdata = 32'd56190;
			9347: outdata = 32'd56189;
			9348: outdata = 32'd56188;
			9349: outdata = 32'd56187;
			9350: outdata = 32'd56186;
			9351: outdata = 32'd56185;
			9352: outdata = 32'd56184;
			9353: outdata = 32'd56183;
			9354: outdata = 32'd56182;
			9355: outdata = 32'd56181;
			9356: outdata = 32'd56180;
			9357: outdata = 32'd56179;
			9358: outdata = 32'd56178;
			9359: outdata = 32'd56177;
			9360: outdata = 32'd56176;
			9361: outdata = 32'd56175;
			9362: outdata = 32'd56174;
			9363: outdata = 32'd56173;
			9364: outdata = 32'd56172;
			9365: outdata = 32'd56171;
			9366: outdata = 32'd56170;
			9367: outdata = 32'd56169;
			9368: outdata = 32'd56168;
			9369: outdata = 32'd56167;
			9370: outdata = 32'd56166;
			9371: outdata = 32'd56165;
			9372: outdata = 32'd56164;
			9373: outdata = 32'd56163;
			9374: outdata = 32'd56162;
			9375: outdata = 32'd56161;
			9376: outdata = 32'd56160;
			9377: outdata = 32'd56159;
			9378: outdata = 32'd56158;
			9379: outdata = 32'd56157;
			9380: outdata = 32'd56156;
			9381: outdata = 32'd56155;
			9382: outdata = 32'd56154;
			9383: outdata = 32'd56153;
			9384: outdata = 32'd56152;
			9385: outdata = 32'd56151;
			9386: outdata = 32'd56150;
			9387: outdata = 32'd56149;
			9388: outdata = 32'd56148;
			9389: outdata = 32'd56147;
			9390: outdata = 32'd56146;
			9391: outdata = 32'd56145;
			9392: outdata = 32'd56144;
			9393: outdata = 32'd56143;
			9394: outdata = 32'd56142;
			9395: outdata = 32'd56141;
			9396: outdata = 32'd56140;
			9397: outdata = 32'd56139;
			9398: outdata = 32'd56138;
			9399: outdata = 32'd56137;
			9400: outdata = 32'd56136;
			9401: outdata = 32'd56135;
			9402: outdata = 32'd56134;
			9403: outdata = 32'd56133;
			9404: outdata = 32'd56132;
			9405: outdata = 32'd56131;
			9406: outdata = 32'd56130;
			9407: outdata = 32'd56129;
			9408: outdata = 32'd56128;
			9409: outdata = 32'd56127;
			9410: outdata = 32'd56126;
			9411: outdata = 32'd56125;
			9412: outdata = 32'd56124;
			9413: outdata = 32'd56123;
			9414: outdata = 32'd56122;
			9415: outdata = 32'd56121;
			9416: outdata = 32'd56120;
			9417: outdata = 32'd56119;
			9418: outdata = 32'd56118;
			9419: outdata = 32'd56117;
			9420: outdata = 32'd56116;
			9421: outdata = 32'd56115;
			9422: outdata = 32'd56114;
			9423: outdata = 32'd56113;
			9424: outdata = 32'd56112;
			9425: outdata = 32'd56111;
			9426: outdata = 32'd56110;
			9427: outdata = 32'd56109;
			9428: outdata = 32'd56108;
			9429: outdata = 32'd56107;
			9430: outdata = 32'd56106;
			9431: outdata = 32'd56105;
			9432: outdata = 32'd56104;
			9433: outdata = 32'd56103;
			9434: outdata = 32'd56102;
			9435: outdata = 32'd56101;
			9436: outdata = 32'd56100;
			9437: outdata = 32'd56099;
			9438: outdata = 32'd56098;
			9439: outdata = 32'd56097;
			9440: outdata = 32'd56096;
			9441: outdata = 32'd56095;
			9442: outdata = 32'd56094;
			9443: outdata = 32'd56093;
			9444: outdata = 32'd56092;
			9445: outdata = 32'd56091;
			9446: outdata = 32'd56090;
			9447: outdata = 32'd56089;
			9448: outdata = 32'd56088;
			9449: outdata = 32'd56087;
			9450: outdata = 32'd56086;
			9451: outdata = 32'd56085;
			9452: outdata = 32'd56084;
			9453: outdata = 32'd56083;
			9454: outdata = 32'd56082;
			9455: outdata = 32'd56081;
			9456: outdata = 32'd56080;
			9457: outdata = 32'd56079;
			9458: outdata = 32'd56078;
			9459: outdata = 32'd56077;
			9460: outdata = 32'd56076;
			9461: outdata = 32'd56075;
			9462: outdata = 32'd56074;
			9463: outdata = 32'd56073;
			9464: outdata = 32'd56072;
			9465: outdata = 32'd56071;
			9466: outdata = 32'd56070;
			9467: outdata = 32'd56069;
			9468: outdata = 32'd56068;
			9469: outdata = 32'd56067;
			9470: outdata = 32'd56066;
			9471: outdata = 32'd56065;
			9472: outdata = 32'd56064;
			9473: outdata = 32'd56063;
			9474: outdata = 32'd56062;
			9475: outdata = 32'd56061;
			9476: outdata = 32'd56060;
			9477: outdata = 32'd56059;
			9478: outdata = 32'd56058;
			9479: outdata = 32'd56057;
			9480: outdata = 32'd56056;
			9481: outdata = 32'd56055;
			9482: outdata = 32'd56054;
			9483: outdata = 32'd56053;
			9484: outdata = 32'd56052;
			9485: outdata = 32'd56051;
			9486: outdata = 32'd56050;
			9487: outdata = 32'd56049;
			9488: outdata = 32'd56048;
			9489: outdata = 32'd56047;
			9490: outdata = 32'd56046;
			9491: outdata = 32'd56045;
			9492: outdata = 32'd56044;
			9493: outdata = 32'd56043;
			9494: outdata = 32'd56042;
			9495: outdata = 32'd56041;
			9496: outdata = 32'd56040;
			9497: outdata = 32'd56039;
			9498: outdata = 32'd56038;
			9499: outdata = 32'd56037;
			9500: outdata = 32'd56036;
			9501: outdata = 32'd56035;
			9502: outdata = 32'd56034;
			9503: outdata = 32'd56033;
			9504: outdata = 32'd56032;
			9505: outdata = 32'd56031;
			9506: outdata = 32'd56030;
			9507: outdata = 32'd56029;
			9508: outdata = 32'd56028;
			9509: outdata = 32'd56027;
			9510: outdata = 32'd56026;
			9511: outdata = 32'd56025;
			9512: outdata = 32'd56024;
			9513: outdata = 32'd56023;
			9514: outdata = 32'd56022;
			9515: outdata = 32'd56021;
			9516: outdata = 32'd56020;
			9517: outdata = 32'd56019;
			9518: outdata = 32'd56018;
			9519: outdata = 32'd56017;
			9520: outdata = 32'd56016;
			9521: outdata = 32'd56015;
			9522: outdata = 32'd56014;
			9523: outdata = 32'd56013;
			9524: outdata = 32'd56012;
			9525: outdata = 32'd56011;
			9526: outdata = 32'd56010;
			9527: outdata = 32'd56009;
			9528: outdata = 32'd56008;
			9529: outdata = 32'd56007;
			9530: outdata = 32'd56006;
			9531: outdata = 32'd56005;
			9532: outdata = 32'd56004;
			9533: outdata = 32'd56003;
			9534: outdata = 32'd56002;
			9535: outdata = 32'd56001;
			9536: outdata = 32'd56000;
			9537: outdata = 32'd55999;
			9538: outdata = 32'd55998;
			9539: outdata = 32'd55997;
			9540: outdata = 32'd55996;
			9541: outdata = 32'd55995;
			9542: outdata = 32'd55994;
			9543: outdata = 32'd55993;
			9544: outdata = 32'd55992;
			9545: outdata = 32'd55991;
			9546: outdata = 32'd55990;
			9547: outdata = 32'd55989;
			9548: outdata = 32'd55988;
			9549: outdata = 32'd55987;
			9550: outdata = 32'd55986;
			9551: outdata = 32'd55985;
			9552: outdata = 32'd55984;
			9553: outdata = 32'd55983;
			9554: outdata = 32'd55982;
			9555: outdata = 32'd55981;
			9556: outdata = 32'd55980;
			9557: outdata = 32'd55979;
			9558: outdata = 32'd55978;
			9559: outdata = 32'd55977;
			9560: outdata = 32'd55976;
			9561: outdata = 32'd55975;
			9562: outdata = 32'd55974;
			9563: outdata = 32'd55973;
			9564: outdata = 32'd55972;
			9565: outdata = 32'd55971;
			9566: outdata = 32'd55970;
			9567: outdata = 32'd55969;
			9568: outdata = 32'd55968;
			9569: outdata = 32'd55967;
			9570: outdata = 32'd55966;
			9571: outdata = 32'd55965;
			9572: outdata = 32'd55964;
			9573: outdata = 32'd55963;
			9574: outdata = 32'd55962;
			9575: outdata = 32'd55961;
			9576: outdata = 32'd55960;
			9577: outdata = 32'd55959;
			9578: outdata = 32'd55958;
			9579: outdata = 32'd55957;
			9580: outdata = 32'd55956;
			9581: outdata = 32'd55955;
			9582: outdata = 32'd55954;
			9583: outdata = 32'd55953;
			9584: outdata = 32'd55952;
			9585: outdata = 32'd55951;
			9586: outdata = 32'd55950;
			9587: outdata = 32'd55949;
			9588: outdata = 32'd55948;
			9589: outdata = 32'd55947;
			9590: outdata = 32'd55946;
			9591: outdata = 32'd55945;
			9592: outdata = 32'd55944;
			9593: outdata = 32'd55943;
			9594: outdata = 32'd55942;
			9595: outdata = 32'd55941;
			9596: outdata = 32'd55940;
			9597: outdata = 32'd55939;
			9598: outdata = 32'd55938;
			9599: outdata = 32'd55937;
			9600: outdata = 32'd55936;
			9601: outdata = 32'd55935;
			9602: outdata = 32'd55934;
			9603: outdata = 32'd55933;
			9604: outdata = 32'd55932;
			9605: outdata = 32'd55931;
			9606: outdata = 32'd55930;
			9607: outdata = 32'd55929;
			9608: outdata = 32'd55928;
			9609: outdata = 32'd55927;
			9610: outdata = 32'd55926;
			9611: outdata = 32'd55925;
			9612: outdata = 32'd55924;
			9613: outdata = 32'd55923;
			9614: outdata = 32'd55922;
			9615: outdata = 32'd55921;
			9616: outdata = 32'd55920;
			9617: outdata = 32'd55919;
			9618: outdata = 32'd55918;
			9619: outdata = 32'd55917;
			9620: outdata = 32'd55916;
			9621: outdata = 32'd55915;
			9622: outdata = 32'd55914;
			9623: outdata = 32'd55913;
			9624: outdata = 32'd55912;
			9625: outdata = 32'd55911;
			9626: outdata = 32'd55910;
			9627: outdata = 32'd55909;
			9628: outdata = 32'd55908;
			9629: outdata = 32'd55907;
			9630: outdata = 32'd55906;
			9631: outdata = 32'd55905;
			9632: outdata = 32'd55904;
			9633: outdata = 32'd55903;
			9634: outdata = 32'd55902;
			9635: outdata = 32'd55901;
			9636: outdata = 32'd55900;
			9637: outdata = 32'd55899;
			9638: outdata = 32'd55898;
			9639: outdata = 32'd55897;
			9640: outdata = 32'd55896;
			9641: outdata = 32'd55895;
			9642: outdata = 32'd55894;
			9643: outdata = 32'd55893;
			9644: outdata = 32'd55892;
			9645: outdata = 32'd55891;
			9646: outdata = 32'd55890;
			9647: outdata = 32'd55889;
			9648: outdata = 32'd55888;
			9649: outdata = 32'd55887;
			9650: outdata = 32'd55886;
			9651: outdata = 32'd55885;
			9652: outdata = 32'd55884;
			9653: outdata = 32'd55883;
			9654: outdata = 32'd55882;
			9655: outdata = 32'd55881;
			9656: outdata = 32'd55880;
			9657: outdata = 32'd55879;
			9658: outdata = 32'd55878;
			9659: outdata = 32'd55877;
			9660: outdata = 32'd55876;
			9661: outdata = 32'd55875;
			9662: outdata = 32'd55874;
			9663: outdata = 32'd55873;
			9664: outdata = 32'd55872;
			9665: outdata = 32'd55871;
			9666: outdata = 32'd55870;
			9667: outdata = 32'd55869;
			9668: outdata = 32'd55868;
			9669: outdata = 32'd55867;
			9670: outdata = 32'd55866;
			9671: outdata = 32'd55865;
			9672: outdata = 32'd55864;
			9673: outdata = 32'd55863;
			9674: outdata = 32'd55862;
			9675: outdata = 32'd55861;
			9676: outdata = 32'd55860;
			9677: outdata = 32'd55859;
			9678: outdata = 32'd55858;
			9679: outdata = 32'd55857;
			9680: outdata = 32'd55856;
			9681: outdata = 32'd55855;
			9682: outdata = 32'd55854;
			9683: outdata = 32'd55853;
			9684: outdata = 32'd55852;
			9685: outdata = 32'd55851;
			9686: outdata = 32'd55850;
			9687: outdata = 32'd55849;
			9688: outdata = 32'd55848;
			9689: outdata = 32'd55847;
			9690: outdata = 32'd55846;
			9691: outdata = 32'd55845;
			9692: outdata = 32'd55844;
			9693: outdata = 32'd55843;
			9694: outdata = 32'd55842;
			9695: outdata = 32'd55841;
			9696: outdata = 32'd55840;
			9697: outdata = 32'd55839;
			9698: outdata = 32'd55838;
			9699: outdata = 32'd55837;
			9700: outdata = 32'd55836;
			9701: outdata = 32'd55835;
			9702: outdata = 32'd55834;
			9703: outdata = 32'd55833;
			9704: outdata = 32'd55832;
			9705: outdata = 32'd55831;
			9706: outdata = 32'd55830;
			9707: outdata = 32'd55829;
			9708: outdata = 32'd55828;
			9709: outdata = 32'd55827;
			9710: outdata = 32'd55826;
			9711: outdata = 32'd55825;
			9712: outdata = 32'd55824;
			9713: outdata = 32'd55823;
			9714: outdata = 32'd55822;
			9715: outdata = 32'd55821;
			9716: outdata = 32'd55820;
			9717: outdata = 32'd55819;
			9718: outdata = 32'd55818;
			9719: outdata = 32'd55817;
			9720: outdata = 32'd55816;
			9721: outdata = 32'd55815;
			9722: outdata = 32'd55814;
			9723: outdata = 32'd55813;
			9724: outdata = 32'd55812;
			9725: outdata = 32'd55811;
			9726: outdata = 32'd55810;
			9727: outdata = 32'd55809;
			9728: outdata = 32'd55808;
			9729: outdata = 32'd55807;
			9730: outdata = 32'd55806;
			9731: outdata = 32'd55805;
			9732: outdata = 32'd55804;
			9733: outdata = 32'd55803;
			9734: outdata = 32'd55802;
			9735: outdata = 32'd55801;
			9736: outdata = 32'd55800;
			9737: outdata = 32'd55799;
			9738: outdata = 32'd55798;
			9739: outdata = 32'd55797;
			9740: outdata = 32'd55796;
			9741: outdata = 32'd55795;
			9742: outdata = 32'd55794;
			9743: outdata = 32'd55793;
			9744: outdata = 32'd55792;
			9745: outdata = 32'd55791;
			9746: outdata = 32'd55790;
			9747: outdata = 32'd55789;
			9748: outdata = 32'd55788;
			9749: outdata = 32'd55787;
			9750: outdata = 32'd55786;
			9751: outdata = 32'd55785;
			9752: outdata = 32'd55784;
			9753: outdata = 32'd55783;
			9754: outdata = 32'd55782;
			9755: outdata = 32'd55781;
			9756: outdata = 32'd55780;
			9757: outdata = 32'd55779;
			9758: outdata = 32'd55778;
			9759: outdata = 32'd55777;
			9760: outdata = 32'd55776;
			9761: outdata = 32'd55775;
			9762: outdata = 32'd55774;
			9763: outdata = 32'd55773;
			9764: outdata = 32'd55772;
			9765: outdata = 32'd55771;
			9766: outdata = 32'd55770;
			9767: outdata = 32'd55769;
			9768: outdata = 32'd55768;
			9769: outdata = 32'd55767;
			9770: outdata = 32'd55766;
			9771: outdata = 32'd55765;
			9772: outdata = 32'd55764;
			9773: outdata = 32'd55763;
			9774: outdata = 32'd55762;
			9775: outdata = 32'd55761;
			9776: outdata = 32'd55760;
			9777: outdata = 32'd55759;
			9778: outdata = 32'd55758;
			9779: outdata = 32'd55757;
			9780: outdata = 32'd55756;
			9781: outdata = 32'd55755;
			9782: outdata = 32'd55754;
			9783: outdata = 32'd55753;
			9784: outdata = 32'd55752;
			9785: outdata = 32'd55751;
			9786: outdata = 32'd55750;
			9787: outdata = 32'd55749;
			9788: outdata = 32'd55748;
			9789: outdata = 32'd55747;
			9790: outdata = 32'd55746;
			9791: outdata = 32'd55745;
			9792: outdata = 32'd55744;
			9793: outdata = 32'd55743;
			9794: outdata = 32'd55742;
			9795: outdata = 32'd55741;
			9796: outdata = 32'd55740;
			9797: outdata = 32'd55739;
			9798: outdata = 32'd55738;
			9799: outdata = 32'd55737;
			9800: outdata = 32'd55736;
			9801: outdata = 32'd55735;
			9802: outdata = 32'd55734;
			9803: outdata = 32'd55733;
			9804: outdata = 32'd55732;
			9805: outdata = 32'd55731;
			9806: outdata = 32'd55730;
			9807: outdata = 32'd55729;
			9808: outdata = 32'd55728;
			9809: outdata = 32'd55727;
			9810: outdata = 32'd55726;
			9811: outdata = 32'd55725;
			9812: outdata = 32'd55724;
			9813: outdata = 32'd55723;
			9814: outdata = 32'd55722;
			9815: outdata = 32'd55721;
			9816: outdata = 32'd55720;
			9817: outdata = 32'd55719;
			9818: outdata = 32'd55718;
			9819: outdata = 32'd55717;
			9820: outdata = 32'd55716;
			9821: outdata = 32'd55715;
			9822: outdata = 32'd55714;
			9823: outdata = 32'd55713;
			9824: outdata = 32'd55712;
			9825: outdata = 32'd55711;
			9826: outdata = 32'd55710;
			9827: outdata = 32'd55709;
			9828: outdata = 32'd55708;
			9829: outdata = 32'd55707;
			9830: outdata = 32'd55706;
			9831: outdata = 32'd55705;
			9832: outdata = 32'd55704;
			9833: outdata = 32'd55703;
			9834: outdata = 32'd55702;
			9835: outdata = 32'd55701;
			9836: outdata = 32'd55700;
			9837: outdata = 32'd55699;
			9838: outdata = 32'd55698;
			9839: outdata = 32'd55697;
			9840: outdata = 32'd55696;
			9841: outdata = 32'd55695;
			9842: outdata = 32'd55694;
			9843: outdata = 32'd55693;
			9844: outdata = 32'd55692;
			9845: outdata = 32'd55691;
			9846: outdata = 32'd55690;
			9847: outdata = 32'd55689;
			9848: outdata = 32'd55688;
			9849: outdata = 32'd55687;
			9850: outdata = 32'd55686;
			9851: outdata = 32'd55685;
			9852: outdata = 32'd55684;
			9853: outdata = 32'd55683;
			9854: outdata = 32'd55682;
			9855: outdata = 32'd55681;
			9856: outdata = 32'd55680;
			9857: outdata = 32'd55679;
			9858: outdata = 32'd55678;
			9859: outdata = 32'd55677;
			9860: outdata = 32'd55676;
			9861: outdata = 32'd55675;
			9862: outdata = 32'd55674;
			9863: outdata = 32'd55673;
			9864: outdata = 32'd55672;
			9865: outdata = 32'd55671;
			9866: outdata = 32'd55670;
			9867: outdata = 32'd55669;
			9868: outdata = 32'd55668;
			9869: outdata = 32'd55667;
			9870: outdata = 32'd55666;
			9871: outdata = 32'd55665;
			9872: outdata = 32'd55664;
			9873: outdata = 32'd55663;
			9874: outdata = 32'd55662;
			9875: outdata = 32'd55661;
			9876: outdata = 32'd55660;
			9877: outdata = 32'd55659;
			9878: outdata = 32'd55658;
			9879: outdata = 32'd55657;
			9880: outdata = 32'd55656;
			9881: outdata = 32'd55655;
			9882: outdata = 32'd55654;
			9883: outdata = 32'd55653;
			9884: outdata = 32'd55652;
			9885: outdata = 32'd55651;
			9886: outdata = 32'd55650;
			9887: outdata = 32'd55649;
			9888: outdata = 32'd55648;
			9889: outdata = 32'd55647;
			9890: outdata = 32'd55646;
			9891: outdata = 32'd55645;
			9892: outdata = 32'd55644;
			9893: outdata = 32'd55643;
			9894: outdata = 32'd55642;
			9895: outdata = 32'd55641;
			9896: outdata = 32'd55640;
			9897: outdata = 32'd55639;
			9898: outdata = 32'd55638;
			9899: outdata = 32'd55637;
			9900: outdata = 32'd55636;
			9901: outdata = 32'd55635;
			9902: outdata = 32'd55634;
			9903: outdata = 32'd55633;
			9904: outdata = 32'd55632;
			9905: outdata = 32'd55631;
			9906: outdata = 32'd55630;
			9907: outdata = 32'd55629;
			9908: outdata = 32'd55628;
			9909: outdata = 32'd55627;
			9910: outdata = 32'd55626;
			9911: outdata = 32'd55625;
			9912: outdata = 32'd55624;
			9913: outdata = 32'd55623;
			9914: outdata = 32'd55622;
			9915: outdata = 32'd55621;
			9916: outdata = 32'd55620;
			9917: outdata = 32'd55619;
			9918: outdata = 32'd55618;
			9919: outdata = 32'd55617;
			9920: outdata = 32'd55616;
			9921: outdata = 32'd55615;
			9922: outdata = 32'd55614;
			9923: outdata = 32'd55613;
			9924: outdata = 32'd55612;
			9925: outdata = 32'd55611;
			9926: outdata = 32'd55610;
			9927: outdata = 32'd55609;
			9928: outdata = 32'd55608;
			9929: outdata = 32'd55607;
			9930: outdata = 32'd55606;
			9931: outdata = 32'd55605;
			9932: outdata = 32'd55604;
			9933: outdata = 32'd55603;
			9934: outdata = 32'd55602;
			9935: outdata = 32'd55601;
			9936: outdata = 32'd55600;
			9937: outdata = 32'd55599;
			9938: outdata = 32'd55598;
			9939: outdata = 32'd55597;
			9940: outdata = 32'd55596;
			9941: outdata = 32'd55595;
			9942: outdata = 32'd55594;
			9943: outdata = 32'd55593;
			9944: outdata = 32'd55592;
			9945: outdata = 32'd55591;
			9946: outdata = 32'd55590;
			9947: outdata = 32'd55589;
			9948: outdata = 32'd55588;
			9949: outdata = 32'd55587;
			9950: outdata = 32'd55586;
			9951: outdata = 32'd55585;
			9952: outdata = 32'd55584;
			9953: outdata = 32'd55583;
			9954: outdata = 32'd55582;
			9955: outdata = 32'd55581;
			9956: outdata = 32'd55580;
			9957: outdata = 32'd55579;
			9958: outdata = 32'd55578;
			9959: outdata = 32'd55577;
			9960: outdata = 32'd55576;
			9961: outdata = 32'd55575;
			9962: outdata = 32'd55574;
			9963: outdata = 32'd55573;
			9964: outdata = 32'd55572;
			9965: outdata = 32'd55571;
			9966: outdata = 32'd55570;
			9967: outdata = 32'd55569;
			9968: outdata = 32'd55568;
			9969: outdata = 32'd55567;
			9970: outdata = 32'd55566;
			9971: outdata = 32'd55565;
			9972: outdata = 32'd55564;
			9973: outdata = 32'd55563;
			9974: outdata = 32'd55562;
			9975: outdata = 32'd55561;
			9976: outdata = 32'd55560;
			9977: outdata = 32'd55559;
			9978: outdata = 32'd55558;
			9979: outdata = 32'd55557;
			9980: outdata = 32'd55556;
			9981: outdata = 32'd55555;
			9982: outdata = 32'd55554;
			9983: outdata = 32'd55553;
			9984: outdata = 32'd55552;
			9985: outdata = 32'd55551;
			9986: outdata = 32'd55550;
			9987: outdata = 32'd55549;
			9988: outdata = 32'd55548;
			9989: outdata = 32'd55547;
			9990: outdata = 32'd55546;
			9991: outdata = 32'd55545;
			9992: outdata = 32'd55544;
			9993: outdata = 32'd55543;
			9994: outdata = 32'd55542;
			9995: outdata = 32'd55541;
			9996: outdata = 32'd55540;
			9997: outdata = 32'd55539;
			9998: outdata = 32'd55538;
			9999: outdata = 32'd55537;
			10000: outdata = 32'd55536;
			10001: outdata = 32'd55535;
			10002: outdata = 32'd55534;
			10003: outdata = 32'd55533;
			10004: outdata = 32'd55532;
			10005: outdata = 32'd55531;
			10006: outdata = 32'd55530;
			10007: outdata = 32'd55529;
			10008: outdata = 32'd55528;
			10009: outdata = 32'd55527;
			10010: outdata = 32'd55526;
			10011: outdata = 32'd55525;
			10012: outdata = 32'd55524;
			10013: outdata = 32'd55523;
			10014: outdata = 32'd55522;
			10015: outdata = 32'd55521;
			10016: outdata = 32'd55520;
			10017: outdata = 32'd55519;
			10018: outdata = 32'd55518;
			10019: outdata = 32'd55517;
			10020: outdata = 32'd55516;
			10021: outdata = 32'd55515;
			10022: outdata = 32'd55514;
			10023: outdata = 32'd55513;
			10024: outdata = 32'd55512;
			10025: outdata = 32'd55511;
			10026: outdata = 32'd55510;
			10027: outdata = 32'd55509;
			10028: outdata = 32'd55508;
			10029: outdata = 32'd55507;
			10030: outdata = 32'd55506;
			10031: outdata = 32'd55505;
			10032: outdata = 32'd55504;
			10033: outdata = 32'd55503;
			10034: outdata = 32'd55502;
			10035: outdata = 32'd55501;
			10036: outdata = 32'd55500;
			10037: outdata = 32'd55499;
			10038: outdata = 32'd55498;
			10039: outdata = 32'd55497;
			10040: outdata = 32'd55496;
			10041: outdata = 32'd55495;
			10042: outdata = 32'd55494;
			10043: outdata = 32'd55493;
			10044: outdata = 32'd55492;
			10045: outdata = 32'd55491;
			10046: outdata = 32'd55490;
			10047: outdata = 32'd55489;
			10048: outdata = 32'd55488;
			10049: outdata = 32'd55487;
			10050: outdata = 32'd55486;
			10051: outdata = 32'd55485;
			10052: outdata = 32'd55484;
			10053: outdata = 32'd55483;
			10054: outdata = 32'd55482;
			10055: outdata = 32'd55481;
			10056: outdata = 32'd55480;
			10057: outdata = 32'd55479;
			10058: outdata = 32'd55478;
			10059: outdata = 32'd55477;
			10060: outdata = 32'd55476;
			10061: outdata = 32'd55475;
			10062: outdata = 32'd55474;
			10063: outdata = 32'd55473;
			10064: outdata = 32'd55472;
			10065: outdata = 32'd55471;
			10066: outdata = 32'd55470;
			10067: outdata = 32'd55469;
			10068: outdata = 32'd55468;
			10069: outdata = 32'd55467;
			10070: outdata = 32'd55466;
			10071: outdata = 32'd55465;
			10072: outdata = 32'd55464;
			10073: outdata = 32'd55463;
			10074: outdata = 32'd55462;
			10075: outdata = 32'd55461;
			10076: outdata = 32'd55460;
			10077: outdata = 32'd55459;
			10078: outdata = 32'd55458;
			10079: outdata = 32'd55457;
			10080: outdata = 32'd55456;
			10081: outdata = 32'd55455;
			10082: outdata = 32'd55454;
			10083: outdata = 32'd55453;
			10084: outdata = 32'd55452;
			10085: outdata = 32'd55451;
			10086: outdata = 32'd55450;
			10087: outdata = 32'd55449;
			10088: outdata = 32'd55448;
			10089: outdata = 32'd55447;
			10090: outdata = 32'd55446;
			10091: outdata = 32'd55445;
			10092: outdata = 32'd55444;
			10093: outdata = 32'd55443;
			10094: outdata = 32'd55442;
			10095: outdata = 32'd55441;
			10096: outdata = 32'd55440;
			10097: outdata = 32'd55439;
			10098: outdata = 32'd55438;
			10099: outdata = 32'd55437;
			10100: outdata = 32'd55436;
			10101: outdata = 32'd55435;
			10102: outdata = 32'd55434;
			10103: outdata = 32'd55433;
			10104: outdata = 32'd55432;
			10105: outdata = 32'd55431;
			10106: outdata = 32'd55430;
			10107: outdata = 32'd55429;
			10108: outdata = 32'd55428;
			10109: outdata = 32'd55427;
			10110: outdata = 32'd55426;
			10111: outdata = 32'd55425;
			10112: outdata = 32'd55424;
			10113: outdata = 32'd55423;
			10114: outdata = 32'd55422;
			10115: outdata = 32'd55421;
			10116: outdata = 32'd55420;
			10117: outdata = 32'd55419;
			10118: outdata = 32'd55418;
			10119: outdata = 32'd55417;
			10120: outdata = 32'd55416;
			10121: outdata = 32'd55415;
			10122: outdata = 32'd55414;
			10123: outdata = 32'd55413;
			10124: outdata = 32'd55412;
			10125: outdata = 32'd55411;
			10126: outdata = 32'd55410;
			10127: outdata = 32'd55409;
			10128: outdata = 32'd55408;
			10129: outdata = 32'd55407;
			10130: outdata = 32'd55406;
			10131: outdata = 32'd55405;
			10132: outdata = 32'd55404;
			10133: outdata = 32'd55403;
			10134: outdata = 32'd55402;
			10135: outdata = 32'd55401;
			10136: outdata = 32'd55400;
			10137: outdata = 32'd55399;
			10138: outdata = 32'd55398;
			10139: outdata = 32'd55397;
			10140: outdata = 32'd55396;
			10141: outdata = 32'd55395;
			10142: outdata = 32'd55394;
			10143: outdata = 32'd55393;
			10144: outdata = 32'd55392;
			10145: outdata = 32'd55391;
			10146: outdata = 32'd55390;
			10147: outdata = 32'd55389;
			10148: outdata = 32'd55388;
			10149: outdata = 32'd55387;
			10150: outdata = 32'd55386;
			10151: outdata = 32'd55385;
			10152: outdata = 32'd55384;
			10153: outdata = 32'd55383;
			10154: outdata = 32'd55382;
			10155: outdata = 32'd55381;
			10156: outdata = 32'd55380;
			10157: outdata = 32'd55379;
			10158: outdata = 32'd55378;
			10159: outdata = 32'd55377;
			10160: outdata = 32'd55376;
			10161: outdata = 32'd55375;
			10162: outdata = 32'd55374;
			10163: outdata = 32'd55373;
			10164: outdata = 32'd55372;
			10165: outdata = 32'd55371;
			10166: outdata = 32'd55370;
			10167: outdata = 32'd55369;
			10168: outdata = 32'd55368;
			10169: outdata = 32'd55367;
			10170: outdata = 32'd55366;
			10171: outdata = 32'd55365;
			10172: outdata = 32'd55364;
			10173: outdata = 32'd55363;
			10174: outdata = 32'd55362;
			10175: outdata = 32'd55361;
			10176: outdata = 32'd55360;
			10177: outdata = 32'd55359;
			10178: outdata = 32'd55358;
			10179: outdata = 32'd55357;
			10180: outdata = 32'd55356;
			10181: outdata = 32'd55355;
			10182: outdata = 32'd55354;
			10183: outdata = 32'd55353;
			10184: outdata = 32'd55352;
			10185: outdata = 32'd55351;
			10186: outdata = 32'd55350;
			10187: outdata = 32'd55349;
			10188: outdata = 32'd55348;
			10189: outdata = 32'd55347;
			10190: outdata = 32'd55346;
			10191: outdata = 32'd55345;
			10192: outdata = 32'd55344;
			10193: outdata = 32'd55343;
			10194: outdata = 32'd55342;
			10195: outdata = 32'd55341;
			10196: outdata = 32'd55340;
			10197: outdata = 32'd55339;
			10198: outdata = 32'd55338;
			10199: outdata = 32'd55337;
			10200: outdata = 32'd55336;
			10201: outdata = 32'd55335;
			10202: outdata = 32'd55334;
			10203: outdata = 32'd55333;
			10204: outdata = 32'd55332;
			10205: outdata = 32'd55331;
			10206: outdata = 32'd55330;
			10207: outdata = 32'd55329;
			10208: outdata = 32'd55328;
			10209: outdata = 32'd55327;
			10210: outdata = 32'd55326;
			10211: outdata = 32'd55325;
			10212: outdata = 32'd55324;
			10213: outdata = 32'd55323;
			10214: outdata = 32'd55322;
			10215: outdata = 32'd55321;
			10216: outdata = 32'd55320;
			10217: outdata = 32'd55319;
			10218: outdata = 32'd55318;
			10219: outdata = 32'd55317;
			10220: outdata = 32'd55316;
			10221: outdata = 32'd55315;
			10222: outdata = 32'd55314;
			10223: outdata = 32'd55313;
			10224: outdata = 32'd55312;
			10225: outdata = 32'd55311;
			10226: outdata = 32'd55310;
			10227: outdata = 32'd55309;
			10228: outdata = 32'd55308;
			10229: outdata = 32'd55307;
			10230: outdata = 32'd55306;
			10231: outdata = 32'd55305;
			10232: outdata = 32'd55304;
			10233: outdata = 32'd55303;
			10234: outdata = 32'd55302;
			10235: outdata = 32'd55301;
			10236: outdata = 32'd55300;
			10237: outdata = 32'd55299;
			10238: outdata = 32'd55298;
			10239: outdata = 32'd55297;
			10240: outdata = 32'd55296;
			10241: outdata = 32'd55295;
			10242: outdata = 32'd55294;
			10243: outdata = 32'd55293;
			10244: outdata = 32'd55292;
			10245: outdata = 32'd55291;
			10246: outdata = 32'd55290;
			10247: outdata = 32'd55289;
			10248: outdata = 32'd55288;
			10249: outdata = 32'd55287;
			10250: outdata = 32'd55286;
			10251: outdata = 32'd55285;
			10252: outdata = 32'd55284;
			10253: outdata = 32'd55283;
			10254: outdata = 32'd55282;
			10255: outdata = 32'd55281;
			10256: outdata = 32'd55280;
			10257: outdata = 32'd55279;
			10258: outdata = 32'd55278;
			10259: outdata = 32'd55277;
			10260: outdata = 32'd55276;
			10261: outdata = 32'd55275;
			10262: outdata = 32'd55274;
			10263: outdata = 32'd55273;
			10264: outdata = 32'd55272;
			10265: outdata = 32'd55271;
			10266: outdata = 32'd55270;
			10267: outdata = 32'd55269;
			10268: outdata = 32'd55268;
			10269: outdata = 32'd55267;
			10270: outdata = 32'd55266;
			10271: outdata = 32'd55265;
			10272: outdata = 32'd55264;
			10273: outdata = 32'd55263;
			10274: outdata = 32'd55262;
			10275: outdata = 32'd55261;
			10276: outdata = 32'd55260;
			10277: outdata = 32'd55259;
			10278: outdata = 32'd55258;
			10279: outdata = 32'd55257;
			10280: outdata = 32'd55256;
			10281: outdata = 32'd55255;
			10282: outdata = 32'd55254;
			10283: outdata = 32'd55253;
			10284: outdata = 32'd55252;
			10285: outdata = 32'd55251;
			10286: outdata = 32'd55250;
			10287: outdata = 32'd55249;
			10288: outdata = 32'd55248;
			10289: outdata = 32'd55247;
			10290: outdata = 32'd55246;
			10291: outdata = 32'd55245;
			10292: outdata = 32'd55244;
			10293: outdata = 32'd55243;
			10294: outdata = 32'd55242;
			10295: outdata = 32'd55241;
			10296: outdata = 32'd55240;
			10297: outdata = 32'd55239;
			10298: outdata = 32'd55238;
			10299: outdata = 32'd55237;
			10300: outdata = 32'd55236;
			10301: outdata = 32'd55235;
			10302: outdata = 32'd55234;
			10303: outdata = 32'd55233;
			10304: outdata = 32'd55232;
			10305: outdata = 32'd55231;
			10306: outdata = 32'd55230;
			10307: outdata = 32'd55229;
			10308: outdata = 32'd55228;
			10309: outdata = 32'd55227;
			10310: outdata = 32'd55226;
			10311: outdata = 32'd55225;
			10312: outdata = 32'd55224;
			10313: outdata = 32'd55223;
			10314: outdata = 32'd55222;
			10315: outdata = 32'd55221;
			10316: outdata = 32'd55220;
			10317: outdata = 32'd55219;
			10318: outdata = 32'd55218;
			10319: outdata = 32'd55217;
			10320: outdata = 32'd55216;
			10321: outdata = 32'd55215;
			10322: outdata = 32'd55214;
			10323: outdata = 32'd55213;
			10324: outdata = 32'd55212;
			10325: outdata = 32'd55211;
			10326: outdata = 32'd55210;
			10327: outdata = 32'd55209;
			10328: outdata = 32'd55208;
			10329: outdata = 32'd55207;
			10330: outdata = 32'd55206;
			10331: outdata = 32'd55205;
			10332: outdata = 32'd55204;
			10333: outdata = 32'd55203;
			10334: outdata = 32'd55202;
			10335: outdata = 32'd55201;
			10336: outdata = 32'd55200;
			10337: outdata = 32'd55199;
			10338: outdata = 32'd55198;
			10339: outdata = 32'd55197;
			10340: outdata = 32'd55196;
			10341: outdata = 32'd55195;
			10342: outdata = 32'd55194;
			10343: outdata = 32'd55193;
			10344: outdata = 32'd55192;
			10345: outdata = 32'd55191;
			10346: outdata = 32'd55190;
			10347: outdata = 32'd55189;
			10348: outdata = 32'd55188;
			10349: outdata = 32'd55187;
			10350: outdata = 32'd55186;
			10351: outdata = 32'd55185;
			10352: outdata = 32'd55184;
			10353: outdata = 32'd55183;
			10354: outdata = 32'd55182;
			10355: outdata = 32'd55181;
			10356: outdata = 32'd55180;
			10357: outdata = 32'd55179;
			10358: outdata = 32'd55178;
			10359: outdata = 32'd55177;
			10360: outdata = 32'd55176;
			10361: outdata = 32'd55175;
			10362: outdata = 32'd55174;
			10363: outdata = 32'd55173;
			10364: outdata = 32'd55172;
			10365: outdata = 32'd55171;
			10366: outdata = 32'd55170;
			10367: outdata = 32'd55169;
			10368: outdata = 32'd55168;
			10369: outdata = 32'd55167;
			10370: outdata = 32'd55166;
			10371: outdata = 32'd55165;
			10372: outdata = 32'd55164;
			10373: outdata = 32'd55163;
			10374: outdata = 32'd55162;
			10375: outdata = 32'd55161;
			10376: outdata = 32'd55160;
			10377: outdata = 32'd55159;
			10378: outdata = 32'd55158;
			10379: outdata = 32'd55157;
			10380: outdata = 32'd55156;
			10381: outdata = 32'd55155;
			10382: outdata = 32'd55154;
			10383: outdata = 32'd55153;
			10384: outdata = 32'd55152;
			10385: outdata = 32'd55151;
			10386: outdata = 32'd55150;
			10387: outdata = 32'd55149;
			10388: outdata = 32'd55148;
			10389: outdata = 32'd55147;
			10390: outdata = 32'd55146;
			10391: outdata = 32'd55145;
			10392: outdata = 32'd55144;
			10393: outdata = 32'd55143;
			10394: outdata = 32'd55142;
			10395: outdata = 32'd55141;
			10396: outdata = 32'd55140;
			10397: outdata = 32'd55139;
			10398: outdata = 32'd55138;
			10399: outdata = 32'd55137;
			10400: outdata = 32'd55136;
			10401: outdata = 32'd55135;
			10402: outdata = 32'd55134;
			10403: outdata = 32'd55133;
			10404: outdata = 32'd55132;
			10405: outdata = 32'd55131;
			10406: outdata = 32'd55130;
			10407: outdata = 32'd55129;
			10408: outdata = 32'd55128;
			10409: outdata = 32'd55127;
			10410: outdata = 32'd55126;
			10411: outdata = 32'd55125;
			10412: outdata = 32'd55124;
			10413: outdata = 32'd55123;
			10414: outdata = 32'd55122;
			10415: outdata = 32'd55121;
			10416: outdata = 32'd55120;
			10417: outdata = 32'd55119;
			10418: outdata = 32'd55118;
			10419: outdata = 32'd55117;
			10420: outdata = 32'd55116;
			10421: outdata = 32'd55115;
			10422: outdata = 32'd55114;
			10423: outdata = 32'd55113;
			10424: outdata = 32'd55112;
			10425: outdata = 32'd55111;
			10426: outdata = 32'd55110;
			10427: outdata = 32'd55109;
			10428: outdata = 32'd55108;
			10429: outdata = 32'd55107;
			10430: outdata = 32'd55106;
			10431: outdata = 32'd55105;
			10432: outdata = 32'd55104;
			10433: outdata = 32'd55103;
			10434: outdata = 32'd55102;
			10435: outdata = 32'd55101;
			10436: outdata = 32'd55100;
			10437: outdata = 32'd55099;
			10438: outdata = 32'd55098;
			10439: outdata = 32'd55097;
			10440: outdata = 32'd55096;
			10441: outdata = 32'd55095;
			10442: outdata = 32'd55094;
			10443: outdata = 32'd55093;
			10444: outdata = 32'd55092;
			10445: outdata = 32'd55091;
			10446: outdata = 32'd55090;
			10447: outdata = 32'd55089;
			10448: outdata = 32'd55088;
			10449: outdata = 32'd55087;
			10450: outdata = 32'd55086;
			10451: outdata = 32'd55085;
			10452: outdata = 32'd55084;
			10453: outdata = 32'd55083;
			10454: outdata = 32'd55082;
			10455: outdata = 32'd55081;
			10456: outdata = 32'd55080;
			10457: outdata = 32'd55079;
			10458: outdata = 32'd55078;
			10459: outdata = 32'd55077;
			10460: outdata = 32'd55076;
			10461: outdata = 32'd55075;
			10462: outdata = 32'd55074;
			10463: outdata = 32'd55073;
			10464: outdata = 32'd55072;
			10465: outdata = 32'd55071;
			10466: outdata = 32'd55070;
			10467: outdata = 32'd55069;
			10468: outdata = 32'd55068;
			10469: outdata = 32'd55067;
			10470: outdata = 32'd55066;
			10471: outdata = 32'd55065;
			10472: outdata = 32'd55064;
			10473: outdata = 32'd55063;
			10474: outdata = 32'd55062;
			10475: outdata = 32'd55061;
			10476: outdata = 32'd55060;
			10477: outdata = 32'd55059;
			10478: outdata = 32'd55058;
			10479: outdata = 32'd55057;
			10480: outdata = 32'd55056;
			10481: outdata = 32'd55055;
			10482: outdata = 32'd55054;
			10483: outdata = 32'd55053;
			10484: outdata = 32'd55052;
			10485: outdata = 32'd55051;
			10486: outdata = 32'd55050;
			10487: outdata = 32'd55049;
			10488: outdata = 32'd55048;
			10489: outdata = 32'd55047;
			10490: outdata = 32'd55046;
			10491: outdata = 32'd55045;
			10492: outdata = 32'd55044;
			10493: outdata = 32'd55043;
			10494: outdata = 32'd55042;
			10495: outdata = 32'd55041;
			10496: outdata = 32'd55040;
			10497: outdata = 32'd55039;
			10498: outdata = 32'd55038;
			10499: outdata = 32'd55037;
			10500: outdata = 32'd55036;
			10501: outdata = 32'd55035;
			10502: outdata = 32'd55034;
			10503: outdata = 32'd55033;
			10504: outdata = 32'd55032;
			10505: outdata = 32'd55031;
			10506: outdata = 32'd55030;
			10507: outdata = 32'd55029;
			10508: outdata = 32'd55028;
			10509: outdata = 32'd55027;
			10510: outdata = 32'd55026;
			10511: outdata = 32'd55025;
			10512: outdata = 32'd55024;
			10513: outdata = 32'd55023;
			10514: outdata = 32'd55022;
			10515: outdata = 32'd55021;
			10516: outdata = 32'd55020;
			10517: outdata = 32'd55019;
			10518: outdata = 32'd55018;
			10519: outdata = 32'd55017;
			10520: outdata = 32'd55016;
			10521: outdata = 32'd55015;
			10522: outdata = 32'd55014;
			10523: outdata = 32'd55013;
			10524: outdata = 32'd55012;
			10525: outdata = 32'd55011;
			10526: outdata = 32'd55010;
			10527: outdata = 32'd55009;
			10528: outdata = 32'd55008;
			10529: outdata = 32'd55007;
			10530: outdata = 32'd55006;
			10531: outdata = 32'd55005;
			10532: outdata = 32'd55004;
			10533: outdata = 32'd55003;
			10534: outdata = 32'd55002;
			10535: outdata = 32'd55001;
			10536: outdata = 32'd55000;
			10537: outdata = 32'd54999;
			10538: outdata = 32'd54998;
			10539: outdata = 32'd54997;
			10540: outdata = 32'd54996;
			10541: outdata = 32'd54995;
			10542: outdata = 32'd54994;
			10543: outdata = 32'd54993;
			10544: outdata = 32'd54992;
			10545: outdata = 32'd54991;
			10546: outdata = 32'd54990;
			10547: outdata = 32'd54989;
			10548: outdata = 32'd54988;
			10549: outdata = 32'd54987;
			10550: outdata = 32'd54986;
			10551: outdata = 32'd54985;
			10552: outdata = 32'd54984;
			10553: outdata = 32'd54983;
			10554: outdata = 32'd54982;
			10555: outdata = 32'd54981;
			10556: outdata = 32'd54980;
			10557: outdata = 32'd54979;
			10558: outdata = 32'd54978;
			10559: outdata = 32'd54977;
			10560: outdata = 32'd54976;
			10561: outdata = 32'd54975;
			10562: outdata = 32'd54974;
			10563: outdata = 32'd54973;
			10564: outdata = 32'd54972;
			10565: outdata = 32'd54971;
			10566: outdata = 32'd54970;
			10567: outdata = 32'd54969;
			10568: outdata = 32'd54968;
			10569: outdata = 32'd54967;
			10570: outdata = 32'd54966;
			10571: outdata = 32'd54965;
			10572: outdata = 32'd54964;
			10573: outdata = 32'd54963;
			10574: outdata = 32'd54962;
			10575: outdata = 32'd54961;
			10576: outdata = 32'd54960;
			10577: outdata = 32'd54959;
			10578: outdata = 32'd54958;
			10579: outdata = 32'd54957;
			10580: outdata = 32'd54956;
			10581: outdata = 32'd54955;
			10582: outdata = 32'd54954;
			10583: outdata = 32'd54953;
			10584: outdata = 32'd54952;
			10585: outdata = 32'd54951;
			10586: outdata = 32'd54950;
			10587: outdata = 32'd54949;
			10588: outdata = 32'd54948;
			10589: outdata = 32'd54947;
			10590: outdata = 32'd54946;
			10591: outdata = 32'd54945;
			10592: outdata = 32'd54944;
			10593: outdata = 32'd54943;
			10594: outdata = 32'd54942;
			10595: outdata = 32'd54941;
			10596: outdata = 32'd54940;
			10597: outdata = 32'd54939;
			10598: outdata = 32'd54938;
			10599: outdata = 32'd54937;
			10600: outdata = 32'd54936;
			10601: outdata = 32'd54935;
			10602: outdata = 32'd54934;
			10603: outdata = 32'd54933;
			10604: outdata = 32'd54932;
			10605: outdata = 32'd54931;
			10606: outdata = 32'd54930;
			10607: outdata = 32'd54929;
			10608: outdata = 32'd54928;
			10609: outdata = 32'd54927;
			10610: outdata = 32'd54926;
			10611: outdata = 32'd54925;
			10612: outdata = 32'd54924;
			10613: outdata = 32'd54923;
			10614: outdata = 32'd54922;
			10615: outdata = 32'd54921;
			10616: outdata = 32'd54920;
			10617: outdata = 32'd54919;
			10618: outdata = 32'd54918;
			10619: outdata = 32'd54917;
			10620: outdata = 32'd54916;
			10621: outdata = 32'd54915;
			10622: outdata = 32'd54914;
			10623: outdata = 32'd54913;
			10624: outdata = 32'd54912;
			10625: outdata = 32'd54911;
			10626: outdata = 32'd54910;
			10627: outdata = 32'd54909;
			10628: outdata = 32'd54908;
			10629: outdata = 32'd54907;
			10630: outdata = 32'd54906;
			10631: outdata = 32'd54905;
			10632: outdata = 32'd54904;
			10633: outdata = 32'd54903;
			10634: outdata = 32'd54902;
			10635: outdata = 32'd54901;
			10636: outdata = 32'd54900;
			10637: outdata = 32'd54899;
			10638: outdata = 32'd54898;
			10639: outdata = 32'd54897;
			10640: outdata = 32'd54896;
			10641: outdata = 32'd54895;
			10642: outdata = 32'd54894;
			10643: outdata = 32'd54893;
			10644: outdata = 32'd54892;
			10645: outdata = 32'd54891;
			10646: outdata = 32'd54890;
			10647: outdata = 32'd54889;
			10648: outdata = 32'd54888;
			10649: outdata = 32'd54887;
			10650: outdata = 32'd54886;
			10651: outdata = 32'd54885;
			10652: outdata = 32'd54884;
			10653: outdata = 32'd54883;
			10654: outdata = 32'd54882;
			10655: outdata = 32'd54881;
			10656: outdata = 32'd54880;
			10657: outdata = 32'd54879;
			10658: outdata = 32'd54878;
			10659: outdata = 32'd54877;
			10660: outdata = 32'd54876;
			10661: outdata = 32'd54875;
			10662: outdata = 32'd54874;
			10663: outdata = 32'd54873;
			10664: outdata = 32'd54872;
			10665: outdata = 32'd54871;
			10666: outdata = 32'd54870;
			10667: outdata = 32'd54869;
			10668: outdata = 32'd54868;
			10669: outdata = 32'd54867;
			10670: outdata = 32'd54866;
			10671: outdata = 32'd54865;
			10672: outdata = 32'd54864;
			10673: outdata = 32'd54863;
			10674: outdata = 32'd54862;
			10675: outdata = 32'd54861;
			10676: outdata = 32'd54860;
			10677: outdata = 32'd54859;
			10678: outdata = 32'd54858;
			10679: outdata = 32'd54857;
			10680: outdata = 32'd54856;
			10681: outdata = 32'd54855;
			10682: outdata = 32'd54854;
			10683: outdata = 32'd54853;
			10684: outdata = 32'd54852;
			10685: outdata = 32'd54851;
			10686: outdata = 32'd54850;
			10687: outdata = 32'd54849;
			10688: outdata = 32'd54848;
			10689: outdata = 32'd54847;
			10690: outdata = 32'd54846;
			10691: outdata = 32'd54845;
			10692: outdata = 32'd54844;
			10693: outdata = 32'd54843;
			10694: outdata = 32'd54842;
			10695: outdata = 32'd54841;
			10696: outdata = 32'd54840;
			10697: outdata = 32'd54839;
			10698: outdata = 32'd54838;
			10699: outdata = 32'd54837;
			10700: outdata = 32'd54836;
			10701: outdata = 32'd54835;
			10702: outdata = 32'd54834;
			10703: outdata = 32'd54833;
			10704: outdata = 32'd54832;
			10705: outdata = 32'd54831;
			10706: outdata = 32'd54830;
			10707: outdata = 32'd54829;
			10708: outdata = 32'd54828;
			10709: outdata = 32'd54827;
			10710: outdata = 32'd54826;
			10711: outdata = 32'd54825;
			10712: outdata = 32'd54824;
			10713: outdata = 32'd54823;
			10714: outdata = 32'd54822;
			10715: outdata = 32'd54821;
			10716: outdata = 32'd54820;
			10717: outdata = 32'd54819;
			10718: outdata = 32'd54818;
			10719: outdata = 32'd54817;
			10720: outdata = 32'd54816;
			10721: outdata = 32'd54815;
			10722: outdata = 32'd54814;
			10723: outdata = 32'd54813;
			10724: outdata = 32'd54812;
			10725: outdata = 32'd54811;
			10726: outdata = 32'd54810;
			10727: outdata = 32'd54809;
			10728: outdata = 32'd54808;
			10729: outdata = 32'd54807;
			10730: outdata = 32'd54806;
			10731: outdata = 32'd54805;
			10732: outdata = 32'd54804;
			10733: outdata = 32'd54803;
			10734: outdata = 32'd54802;
			10735: outdata = 32'd54801;
			10736: outdata = 32'd54800;
			10737: outdata = 32'd54799;
			10738: outdata = 32'd54798;
			10739: outdata = 32'd54797;
			10740: outdata = 32'd54796;
			10741: outdata = 32'd54795;
			10742: outdata = 32'd54794;
			10743: outdata = 32'd54793;
			10744: outdata = 32'd54792;
			10745: outdata = 32'd54791;
			10746: outdata = 32'd54790;
			10747: outdata = 32'd54789;
			10748: outdata = 32'd54788;
			10749: outdata = 32'd54787;
			10750: outdata = 32'd54786;
			10751: outdata = 32'd54785;
			10752: outdata = 32'd54784;
			10753: outdata = 32'd54783;
			10754: outdata = 32'd54782;
			10755: outdata = 32'd54781;
			10756: outdata = 32'd54780;
			10757: outdata = 32'd54779;
			10758: outdata = 32'd54778;
			10759: outdata = 32'd54777;
			10760: outdata = 32'd54776;
			10761: outdata = 32'd54775;
			10762: outdata = 32'd54774;
			10763: outdata = 32'd54773;
			10764: outdata = 32'd54772;
			10765: outdata = 32'd54771;
			10766: outdata = 32'd54770;
			10767: outdata = 32'd54769;
			10768: outdata = 32'd54768;
			10769: outdata = 32'd54767;
			10770: outdata = 32'd54766;
			10771: outdata = 32'd54765;
			10772: outdata = 32'd54764;
			10773: outdata = 32'd54763;
			10774: outdata = 32'd54762;
			10775: outdata = 32'd54761;
			10776: outdata = 32'd54760;
			10777: outdata = 32'd54759;
			10778: outdata = 32'd54758;
			10779: outdata = 32'd54757;
			10780: outdata = 32'd54756;
			10781: outdata = 32'd54755;
			10782: outdata = 32'd54754;
			10783: outdata = 32'd54753;
			10784: outdata = 32'd54752;
			10785: outdata = 32'd54751;
			10786: outdata = 32'd54750;
			10787: outdata = 32'd54749;
			10788: outdata = 32'd54748;
			10789: outdata = 32'd54747;
			10790: outdata = 32'd54746;
			10791: outdata = 32'd54745;
			10792: outdata = 32'd54744;
			10793: outdata = 32'd54743;
			10794: outdata = 32'd54742;
			10795: outdata = 32'd54741;
			10796: outdata = 32'd54740;
			10797: outdata = 32'd54739;
			10798: outdata = 32'd54738;
			10799: outdata = 32'd54737;
			10800: outdata = 32'd54736;
			10801: outdata = 32'd54735;
			10802: outdata = 32'd54734;
			10803: outdata = 32'd54733;
			10804: outdata = 32'd54732;
			10805: outdata = 32'd54731;
			10806: outdata = 32'd54730;
			10807: outdata = 32'd54729;
			10808: outdata = 32'd54728;
			10809: outdata = 32'd54727;
			10810: outdata = 32'd54726;
			10811: outdata = 32'd54725;
			10812: outdata = 32'd54724;
			10813: outdata = 32'd54723;
			10814: outdata = 32'd54722;
			10815: outdata = 32'd54721;
			10816: outdata = 32'd54720;
			10817: outdata = 32'd54719;
			10818: outdata = 32'd54718;
			10819: outdata = 32'd54717;
			10820: outdata = 32'd54716;
			10821: outdata = 32'd54715;
			10822: outdata = 32'd54714;
			10823: outdata = 32'd54713;
			10824: outdata = 32'd54712;
			10825: outdata = 32'd54711;
			10826: outdata = 32'd54710;
			10827: outdata = 32'd54709;
			10828: outdata = 32'd54708;
			10829: outdata = 32'd54707;
			10830: outdata = 32'd54706;
			10831: outdata = 32'd54705;
			10832: outdata = 32'd54704;
			10833: outdata = 32'd54703;
			10834: outdata = 32'd54702;
			10835: outdata = 32'd54701;
			10836: outdata = 32'd54700;
			10837: outdata = 32'd54699;
			10838: outdata = 32'd54698;
			10839: outdata = 32'd54697;
			10840: outdata = 32'd54696;
			10841: outdata = 32'd54695;
			10842: outdata = 32'd54694;
			10843: outdata = 32'd54693;
			10844: outdata = 32'd54692;
			10845: outdata = 32'd54691;
			10846: outdata = 32'd54690;
			10847: outdata = 32'd54689;
			10848: outdata = 32'd54688;
			10849: outdata = 32'd54687;
			10850: outdata = 32'd54686;
			10851: outdata = 32'd54685;
			10852: outdata = 32'd54684;
			10853: outdata = 32'd54683;
			10854: outdata = 32'd54682;
			10855: outdata = 32'd54681;
			10856: outdata = 32'd54680;
			10857: outdata = 32'd54679;
			10858: outdata = 32'd54678;
			10859: outdata = 32'd54677;
			10860: outdata = 32'd54676;
			10861: outdata = 32'd54675;
			10862: outdata = 32'd54674;
			10863: outdata = 32'd54673;
			10864: outdata = 32'd54672;
			10865: outdata = 32'd54671;
			10866: outdata = 32'd54670;
			10867: outdata = 32'd54669;
			10868: outdata = 32'd54668;
			10869: outdata = 32'd54667;
			10870: outdata = 32'd54666;
			10871: outdata = 32'd54665;
			10872: outdata = 32'd54664;
			10873: outdata = 32'd54663;
			10874: outdata = 32'd54662;
			10875: outdata = 32'd54661;
			10876: outdata = 32'd54660;
			10877: outdata = 32'd54659;
			10878: outdata = 32'd54658;
			10879: outdata = 32'd54657;
			10880: outdata = 32'd54656;
			10881: outdata = 32'd54655;
			10882: outdata = 32'd54654;
			10883: outdata = 32'd54653;
			10884: outdata = 32'd54652;
			10885: outdata = 32'd54651;
			10886: outdata = 32'd54650;
			10887: outdata = 32'd54649;
			10888: outdata = 32'd54648;
			10889: outdata = 32'd54647;
			10890: outdata = 32'd54646;
			10891: outdata = 32'd54645;
			10892: outdata = 32'd54644;
			10893: outdata = 32'd54643;
			10894: outdata = 32'd54642;
			10895: outdata = 32'd54641;
			10896: outdata = 32'd54640;
			10897: outdata = 32'd54639;
			10898: outdata = 32'd54638;
			10899: outdata = 32'd54637;
			10900: outdata = 32'd54636;
			10901: outdata = 32'd54635;
			10902: outdata = 32'd54634;
			10903: outdata = 32'd54633;
			10904: outdata = 32'd54632;
			10905: outdata = 32'd54631;
			10906: outdata = 32'd54630;
			10907: outdata = 32'd54629;
			10908: outdata = 32'd54628;
			10909: outdata = 32'd54627;
			10910: outdata = 32'd54626;
			10911: outdata = 32'd54625;
			10912: outdata = 32'd54624;
			10913: outdata = 32'd54623;
			10914: outdata = 32'd54622;
			10915: outdata = 32'd54621;
			10916: outdata = 32'd54620;
			10917: outdata = 32'd54619;
			10918: outdata = 32'd54618;
			10919: outdata = 32'd54617;
			10920: outdata = 32'd54616;
			10921: outdata = 32'd54615;
			10922: outdata = 32'd54614;
			10923: outdata = 32'd54613;
			10924: outdata = 32'd54612;
			10925: outdata = 32'd54611;
			10926: outdata = 32'd54610;
			10927: outdata = 32'd54609;
			10928: outdata = 32'd54608;
			10929: outdata = 32'd54607;
			10930: outdata = 32'd54606;
			10931: outdata = 32'd54605;
			10932: outdata = 32'd54604;
			10933: outdata = 32'd54603;
			10934: outdata = 32'd54602;
			10935: outdata = 32'd54601;
			10936: outdata = 32'd54600;
			10937: outdata = 32'd54599;
			10938: outdata = 32'd54598;
			10939: outdata = 32'd54597;
			10940: outdata = 32'd54596;
			10941: outdata = 32'd54595;
			10942: outdata = 32'd54594;
			10943: outdata = 32'd54593;
			10944: outdata = 32'd54592;
			10945: outdata = 32'd54591;
			10946: outdata = 32'd54590;
			10947: outdata = 32'd54589;
			10948: outdata = 32'd54588;
			10949: outdata = 32'd54587;
			10950: outdata = 32'd54586;
			10951: outdata = 32'd54585;
			10952: outdata = 32'd54584;
			10953: outdata = 32'd54583;
			10954: outdata = 32'd54582;
			10955: outdata = 32'd54581;
			10956: outdata = 32'd54580;
			10957: outdata = 32'd54579;
			10958: outdata = 32'd54578;
			10959: outdata = 32'd54577;
			10960: outdata = 32'd54576;
			10961: outdata = 32'd54575;
			10962: outdata = 32'd54574;
			10963: outdata = 32'd54573;
			10964: outdata = 32'd54572;
			10965: outdata = 32'd54571;
			10966: outdata = 32'd54570;
			10967: outdata = 32'd54569;
			10968: outdata = 32'd54568;
			10969: outdata = 32'd54567;
			10970: outdata = 32'd54566;
			10971: outdata = 32'd54565;
			10972: outdata = 32'd54564;
			10973: outdata = 32'd54563;
			10974: outdata = 32'd54562;
			10975: outdata = 32'd54561;
			10976: outdata = 32'd54560;
			10977: outdata = 32'd54559;
			10978: outdata = 32'd54558;
			10979: outdata = 32'd54557;
			10980: outdata = 32'd54556;
			10981: outdata = 32'd54555;
			10982: outdata = 32'd54554;
			10983: outdata = 32'd54553;
			10984: outdata = 32'd54552;
			10985: outdata = 32'd54551;
			10986: outdata = 32'd54550;
			10987: outdata = 32'd54549;
			10988: outdata = 32'd54548;
			10989: outdata = 32'd54547;
			10990: outdata = 32'd54546;
			10991: outdata = 32'd54545;
			10992: outdata = 32'd54544;
			10993: outdata = 32'd54543;
			10994: outdata = 32'd54542;
			10995: outdata = 32'd54541;
			10996: outdata = 32'd54540;
			10997: outdata = 32'd54539;
			10998: outdata = 32'd54538;
			10999: outdata = 32'd54537;
			11000: outdata = 32'd54536;
			11001: outdata = 32'd54535;
			11002: outdata = 32'd54534;
			11003: outdata = 32'd54533;
			11004: outdata = 32'd54532;
			11005: outdata = 32'd54531;
			11006: outdata = 32'd54530;
			11007: outdata = 32'd54529;
			11008: outdata = 32'd54528;
			11009: outdata = 32'd54527;
			11010: outdata = 32'd54526;
			11011: outdata = 32'd54525;
			11012: outdata = 32'd54524;
			11013: outdata = 32'd54523;
			11014: outdata = 32'd54522;
			11015: outdata = 32'd54521;
			11016: outdata = 32'd54520;
			11017: outdata = 32'd54519;
			11018: outdata = 32'd54518;
			11019: outdata = 32'd54517;
			11020: outdata = 32'd54516;
			11021: outdata = 32'd54515;
			11022: outdata = 32'd54514;
			11023: outdata = 32'd54513;
			11024: outdata = 32'd54512;
			11025: outdata = 32'd54511;
			11026: outdata = 32'd54510;
			11027: outdata = 32'd54509;
			11028: outdata = 32'd54508;
			11029: outdata = 32'd54507;
			11030: outdata = 32'd54506;
			11031: outdata = 32'd54505;
			11032: outdata = 32'd54504;
			11033: outdata = 32'd54503;
			11034: outdata = 32'd54502;
			11035: outdata = 32'd54501;
			11036: outdata = 32'd54500;
			11037: outdata = 32'd54499;
			11038: outdata = 32'd54498;
			11039: outdata = 32'd54497;
			11040: outdata = 32'd54496;
			11041: outdata = 32'd54495;
			11042: outdata = 32'd54494;
			11043: outdata = 32'd54493;
			11044: outdata = 32'd54492;
			11045: outdata = 32'd54491;
			11046: outdata = 32'd54490;
			11047: outdata = 32'd54489;
			11048: outdata = 32'd54488;
			11049: outdata = 32'd54487;
			11050: outdata = 32'd54486;
			11051: outdata = 32'd54485;
			11052: outdata = 32'd54484;
			11053: outdata = 32'd54483;
			11054: outdata = 32'd54482;
			11055: outdata = 32'd54481;
			11056: outdata = 32'd54480;
			11057: outdata = 32'd54479;
			11058: outdata = 32'd54478;
			11059: outdata = 32'd54477;
			11060: outdata = 32'd54476;
			11061: outdata = 32'd54475;
			11062: outdata = 32'd54474;
			11063: outdata = 32'd54473;
			11064: outdata = 32'd54472;
			11065: outdata = 32'd54471;
			11066: outdata = 32'd54470;
			11067: outdata = 32'd54469;
			11068: outdata = 32'd54468;
			11069: outdata = 32'd54467;
			11070: outdata = 32'd54466;
			11071: outdata = 32'd54465;
			11072: outdata = 32'd54464;
			11073: outdata = 32'd54463;
			11074: outdata = 32'd54462;
			11075: outdata = 32'd54461;
			11076: outdata = 32'd54460;
			11077: outdata = 32'd54459;
			11078: outdata = 32'd54458;
			11079: outdata = 32'd54457;
			11080: outdata = 32'd54456;
			11081: outdata = 32'd54455;
			11082: outdata = 32'd54454;
			11083: outdata = 32'd54453;
			11084: outdata = 32'd54452;
			11085: outdata = 32'd54451;
			11086: outdata = 32'd54450;
			11087: outdata = 32'd54449;
			11088: outdata = 32'd54448;
			11089: outdata = 32'd54447;
			11090: outdata = 32'd54446;
			11091: outdata = 32'd54445;
			11092: outdata = 32'd54444;
			11093: outdata = 32'd54443;
			11094: outdata = 32'd54442;
			11095: outdata = 32'd54441;
			11096: outdata = 32'd54440;
			11097: outdata = 32'd54439;
			11098: outdata = 32'd54438;
			11099: outdata = 32'd54437;
			11100: outdata = 32'd54436;
			11101: outdata = 32'd54435;
			11102: outdata = 32'd54434;
			11103: outdata = 32'd54433;
			11104: outdata = 32'd54432;
			11105: outdata = 32'd54431;
			11106: outdata = 32'd54430;
			11107: outdata = 32'd54429;
			11108: outdata = 32'd54428;
			11109: outdata = 32'd54427;
			11110: outdata = 32'd54426;
			11111: outdata = 32'd54425;
			11112: outdata = 32'd54424;
			11113: outdata = 32'd54423;
			11114: outdata = 32'd54422;
			11115: outdata = 32'd54421;
			11116: outdata = 32'd54420;
			11117: outdata = 32'd54419;
			11118: outdata = 32'd54418;
			11119: outdata = 32'd54417;
			11120: outdata = 32'd54416;
			11121: outdata = 32'd54415;
			11122: outdata = 32'd54414;
			11123: outdata = 32'd54413;
			11124: outdata = 32'd54412;
			11125: outdata = 32'd54411;
			11126: outdata = 32'd54410;
			11127: outdata = 32'd54409;
			11128: outdata = 32'd54408;
			11129: outdata = 32'd54407;
			11130: outdata = 32'd54406;
			11131: outdata = 32'd54405;
			11132: outdata = 32'd54404;
			11133: outdata = 32'd54403;
			11134: outdata = 32'd54402;
			11135: outdata = 32'd54401;
			11136: outdata = 32'd54400;
			11137: outdata = 32'd54399;
			11138: outdata = 32'd54398;
			11139: outdata = 32'd54397;
			11140: outdata = 32'd54396;
			11141: outdata = 32'd54395;
			11142: outdata = 32'd54394;
			11143: outdata = 32'd54393;
			11144: outdata = 32'd54392;
			11145: outdata = 32'd54391;
			11146: outdata = 32'd54390;
			11147: outdata = 32'd54389;
			11148: outdata = 32'd54388;
			11149: outdata = 32'd54387;
			11150: outdata = 32'd54386;
			11151: outdata = 32'd54385;
			11152: outdata = 32'd54384;
			11153: outdata = 32'd54383;
			11154: outdata = 32'd54382;
			11155: outdata = 32'd54381;
			11156: outdata = 32'd54380;
			11157: outdata = 32'd54379;
			11158: outdata = 32'd54378;
			11159: outdata = 32'd54377;
			11160: outdata = 32'd54376;
			11161: outdata = 32'd54375;
			11162: outdata = 32'd54374;
			11163: outdata = 32'd54373;
			11164: outdata = 32'd54372;
			11165: outdata = 32'd54371;
			11166: outdata = 32'd54370;
			11167: outdata = 32'd54369;
			11168: outdata = 32'd54368;
			11169: outdata = 32'd54367;
			11170: outdata = 32'd54366;
			11171: outdata = 32'd54365;
			11172: outdata = 32'd54364;
			11173: outdata = 32'd54363;
			11174: outdata = 32'd54362;
			11175: outdata = 32'd54361;
			11176: outdata = 32'd54360;
			11177: outdata = 32'd54359;
			11178: outdata = 32'd54358;
			11179: outdata = 32'd54357;
			11180: outdata = 32'd54356;
			11181: outdata = 32'd54355;
			11182: outdata = 32'd54354;
			11183: outdata = 32'd54353;
			11184: outdata = 32'd54352;
			11185: outdata = 32'd54351;
			11186: outdata = 32'd54350;
			11187: outdata = 32'd54349;
			11188: outdata = 32'd54348;
			11189: outdata = 32'd54347;
			11190: outdata = 32'd54346;
			11191: outdata = 32'd54345;
			11192: outdata = 32'd54344;
			11193: outdata = 32'd54343;
			11194: outdata = 32'd54342;
			11195: outdata = 32'd54341;
			11196: outdata = 32'd54340;
			11197: outdata = 32'd54339;
			11198: outdata = 32'd54338;
			11199: outdata = 32'd54337;
			11200: outdata = 32'd54336;
			11201: outdata = 32'd54335;
			11202: outdata = 32'd54334;
			11203: outdata = 32'd54333;
			11204: outdata = 32'd54332;
			11205: outdata = 32'd54331;
			11206: outdata = 32'd54330;
			11207: outdata = 32'd54329;
			11208: outdata = 32'd54328;
			11209: outdata = 32'd54327;
			11210: outdata = 32'd54326;
			11211: outdata = 32'd54325;
			11212: outdata = 32'd54324;
			11213: outdata = 32'd54323;
			11214: outdata = 32'd54322;
			11215: outdata = 32'd54321;
			11216: outdata = 32'd54320;
			11217: outdata = 32'd54319;
			11218: outdata = 32'd54318;
			11219: outdata = 32'd54317;
			11220: outdata = 32'd54316;
			11221: outdata = 32'd54315;
			11222: outdata = 32'd54314;
			11223: outdata = 32'd54313;
			11224: outdata = 32'd54312;
			11225: outdata = 32'd54311;
			11226: outdata = 32'd54310;
			11227: outdata = 32'd54309;
			11228: outdata = 32'd54308;
			11229: outdata = 32'd54307;
			11230: outdata = 32'd54306;
			11231: outdata = 32'd54305;
			11232: outdata = 32'd54304;
			11233: outdata = 32'd54303;
			11234: outdata = 32'd54302;
			11235: outdata = 32'd54301;
			11236: outdata = 32'd54300;
			11237: outdata = 32'd54299;
			11238: outdata = 32'd54298;
			11239: outdata = 32'd54297;
			11240: outdata = 32'd54296;
			11241: outdata = 32'd54295;
			11242: outdata = 32'd54294;
			11243: outdata = 32'd54293;
			11244: outdata = 32'd54292;
			11245: outdata = 32'd54291;
			11246: outdata = 32'd54290;
			11247: outdata = 32'd54289;
			11248: outdata = 32'd54288;
			11249: outdata = 32'd54287;
			11250: outdata = 32'd54286;
			11251: outdata = 32'd54285;
			11252: outdata = 32'd54284;
			11253: outdata = 32'd54283;
			11254: outdata = 32'd54282;
			11255: outdata = 32'd54281;
			11256: outdata = 32'd54280;
			11257: outdata = 32'd54279;
			11258: outdata = 32'd54278;
			11259: outdata = 32'd54277;
			11260: outdata = 32'd54276;
			11261: outdata = 32'd54275;
			11262: outdata = 32'd54274;
			11263: outdata = 32'd54273;
			11264: outdata = 32'd54272;
			11265: outdata = 32'd54271;
			11266: outdata = 32'd54270;
			11267: outdata = 32'd54269;
			11268: outdata = 32'd54268;
			11269: outdata = 32'd54267;
			11270: outdata = 32'd54266;
			11271: outdata = 32'd54265;
			11272: outdata = 32'd54264;
			11273: outdata = 32'd54263;
			11274: outdata = 32'd54262;
			11275: outdata = 32'd54261;
			11276: outdata = 32'd54260;
			11277: outdata = 32'd54259;
			11278: outdata = 32'd54258;
			11279: outdata = 32'd54257;
			11280: outdata = 32'd54256;
			11281: outdata = 32'd54255;
			11282: outdata = 32'd54254;
			11283: outdata = 32'd54253;
			11284: outdata = 32'd54252;
			11285: outdata = 32'd54251;
			11286: outdata = 32'd54250;
			11287: outdata = 32'd54249;
			11288: outdata = 32'd54248;
			11289: outdata = 32'd54247;
			11290: outdata = 32'd54246;
			11291: outdata = 32'd54245;
			11292: outdata = 32'd54244;
			11293: outdata = 32'd54243;
			11294: outdata = 32'd54242;
			11295: outdata = 32'd54241;
			11296: outdata = 32'd54240;
			11297: outdata = 32'd54239;
			11298: outdata = 32'd54238;
			11299: outdata = 32'd54237;
			11300: outdata = 32'd54236;
			11301: outdata = 32'd54235;
			11302: outdata = 32'd54234;
			11303: outdata = 32'd54233;
			11304: outdata = 32'd54232;
			11305: outdata = 32'd54231;
			11306: outdata = 32'd54230;
			11307: outdata = 32'd54229;
			11308: outdata = 32'd54228;
			11309: outdata = 32'd54227;
			11310: outdata = 32'd54226;
			11311: outdata = 32'd54225;
			11312: outdata = 32'd54224;
			11313: outdata = 32'd54223;
			11314: outdata = 32'd54222;
			11315: outdata = 32'd54221;
			11316: outdata = 32'd54220;
			11317: outdata = 32'd54219;
			11318: outdata = 32'd54218;
			11319: outdata = 32'd54217;
			11320: outdata = 32'd54216;
			11321: outdata = 32'd54215;
			11322: outdata = 32'd54214;
			11323: outdata = 32'd54213;
			11324: outdata = 32'd54212;
			11325: outdata = 32'd54211;
			11326: outdata = 32'd54210;
			11327: outdata = 32'd54209;
			11328: outdata = 32'd54208;
			11329: outdata = 32'd54207;
			11330: outdata = 32'd54206;
			11331: outdata = 32'd54205;
			11332: outdata = 32'd54204;
			11333: outdata = 32'd54203;
			11334: outdata = 32'd54202;
			11335: outdata = 32'd54201;
			11336: outdata = 32'd54200;
			11337: outdata = 32'd54199;
			11338: outdata = 32'd54198;
			11339: outdata = 32'd54197;
			11340: outdata = 32'd54196;
			11341: outdata = 32'd54195;
			11342: outdata = 32'd54194;
			11343: outdata = 32'd54193;
			11344: outdata = 32'd54192;
			11345: outdata = 32'd54191;
			11346: outdata = 32'd54190;
			11347: outdata = 32'd54189;
			11348: outdata = 32'd54188;
			11349: outdata = 32'd54187;
			11350: outdata = 32'd54186;
			11351: outdata = 32'd54185;
			11352: outdata = 32'd54184;
			11353: outdata = 32'd54183;
			11354: outdata = 32'd54182;
			11355: outdata = 32'd54181;
			11356: outdata = 32'd54180;
			11357: outdata = 32'd54179;
			11358: outdata = 32'd54178;
			11359: outdata = 32'd54177;
			11360: outdata = 32'd54176;
			11361: outdata = 32'd54175;
			11362: outdata = 32'd54174;
			11363: outdata = 32'd54173;
			11364: outdata = 32'd54172;
			11365: outdata = 32'd54171;
			11366: outdata = 32'd54170;
			11367: outdata = 32'd54169;
			11368: outdata = 32'd54168;
			11369: outdata = 32'd54167;
			11370: outdata = 32'd54166;
			11371: outdata = 32'd54165;
			11372: outdata = 32'd54164;
			11373: outdata = 32'd54163;
			11374: outdata = 32'd54162;
			11375: outdata = 32'd54161;
			11376: outdata = 32'd54160;
			11377: outdata = 32'd54159;
			11378: outdata = 32'd54158;
			11379: outdata = 32'd54157;
			11380: outdata = 32'd54156;
			11381: outdata = 32'd54155;
			11382: outdata = 32'd54154;
			11383: outdata = 32'd54153;
			11384: outdata = 32'd54152;
			11385: outdata = 32'd54151;
			11386: outdata = 32'd54150;
			11387: outdata = 32'd54149;
			11388: outdata = 32'd54148;
			11389: outdata = 32'd54147;
			11390: outdata = 32'd54146;
			11391: outdata = 32'd54145;
			11392: outdata = 32'd54144;
			11393: outdata = 32'd54143;
			11394: outdata = 32'd54142;
			11395: outdata = 32'd54141;
			11396: outdata = 32'd54140;
			11397: outdata = 32'd54139;
			11398: outdata = 32'd54138;
			11399: outdata = 32'd54137;
			11400: outdata = 32'd54136;
			11401: outdata = 32'd54135;
			11402: outdata = 32'd54134;
			11403: outdata = 32'd54133;
			11404: outdata = 32'd54132;
			11405: outdata = 32'd54131;
			11406: outdata = 32'd54130;
			11407: outdata = 32'd54129;
			11408: outdata = 32'd54128;
			11409: outdata = 32'd54127;
			11410: outdata = 32'd54126;
			11411: outdata = 32'd54125;
			11412: outdata = 32'd54124;
			11413: outdata = 32'd54123;
			11414: outdata = 32'd54122;
			11415: outdata = 32'd54121;
			11416: outdata = 32'd54120;
			11417: outdata = 32'd54119;
			11418: outdata = 32'd54118;
			11419: outdata = 32'd54117;
			11420: outdata = 32'd54116;
			11421: outdata = 32'd54115;
			11422: outdata = 32'd54114;
			11423: outdata = 32'd54113;
			11424: outdata = 32'd54112;
			11425: outdata = 32'd54111;
			11426: outdata = 32'd54110;
			11427: outdata = 32'd54109;
			11428: outdata = 32'd54108;
			11429: outdata = 32'd54107;
			11430: outdata = 32'd54106;
			11431: outdata = 32'd54105;
			11432: outdata = 32'd54104;
			11433: outdata = 32'd54103;
			11434: outdata = 32'd54102;
			11435: outdata = 32'd54101;
			11436: outdata = 32'd54100;
			11437: outdata = 32'd54099;
			11438: outdata = 32'd54098;
			11439: outdata = 32'd54097;
			11440: outdata = 32'd54096;
			11441: outdata = 32'd54095;
			11442: outdata = 32'd54094;
			11443: outdata = 32'd54093;
			11444: outdata = 32'd54092;
			11445: outdata = 32'd54091;
			11446: outdata = 32'd54090;
			11447: outdata = 32'd54089;
			11448: outdata = 32'd54088;
			11449: outdata = 32'd54087;
			11450: outdata = 32'd54086;
			11451: outdata = 32'd54085;
			11452: outdata = 32'd54084;
			11453: outdata = 32'd54083;
			11454: outdata = 32'd54082;
			11455: outdata = 32'd54081;
			11456: outdata = 32'd54080;
			11457: outdata = 32'd54079;
			11458: outdata = 32'd54078;
			11459: outdata = 32'd54077;
			11460: outdata = 32'd54076;
			11461: outdata = 32'd54075;
			11462: outdata = 32'd54074;
			11463: outdata = 32'd54073;
			11464: outdata = 32'd54072;
			11465: outdata = 32'd54071;
			11466: outdata = 32'd54070;
			11467: outdata = 32'd54069;
			11468: outdata = 32'd54068;
			11469: outdata = 32'd54067;
			11470: outdata = 32'd54066;
			11471: outdata = 32'd54065;
			11472: outdata = 32'd54064;
			11473: outdata = 32'd54063;
			11474: outdata = 32'd54062;
			11475: outdata = 32'd54061;
			11476: outdata = 32'd54060;
			11477: outdata = 32'd54059;
			11478: outdata = 32'd54058;
			11479: outdata = 32'd54057;
			11480: outdata = 32'd54056;
			11481: outdata = 32'd54055;
			11482: outdata = 32'd54054;
			11483: outdata = 32'd54053;
			11484: outdata = 32'd54052;
			11485: outdata = 32'd54051;
			11486: outdata = 32'd54050;
			11487: outdata = 32'd54049;
			11488: outdata = 32'd54048;
			11489: outdata = 32'd54047;
			11490: outdata = 32'd54046;
			11491: outdata = 32'd54045;
			11492: outdata = 32'd54044;
			11493: outdata = 32'd54043;
			11494: outdata = 32'd54042;
			11495: outdata = 32'd54041;
			11496: outdata = 32'd54040;
			11497: outdata = 32'd54039;
			11498: outdata = 32'd54038;
			11499: outdata = 32'd54037;
			11500: outdata = 32'd54036;
			11501: outdata = 32'd54035;
			11502: outdata = 32'd54034;
			11503: outdata = 32'd54033;
			11504: outdata = 32'd54032;
			11505: outdata = 32'd54031;
			11506: outdata = 32'd54030;
			11507: outdata = 32'd54029;
			11508: outdata = 32'd54028;
			11509: outdata = 32'd54027;
			11510: outdata = 32'd54026;
			11511: outdata = 32'd54025;
			11512: outdata = 32'd54024;
			11513: outdata = 32'd54023;
			11514: outdata = 32'd54022;
			11515: outdata = 32'd54021;
			11516: outdata = 32'd54020;
			11517: outdata = 32'd54019;
			11518: outdata = 32'd54018;
			11519: outdata = 32'd54017;
			11520: outdata = 32'd54016;
			11521: outdata = 32'd54015;
			11522: outdata = 32'd54014;
			11523: outdata = 32'd54013;
			11524: outdata = 32'd54012;
			11525: outdata = 32'd54011;
			11526: outdata = 32'd54010;
			11527: outdata = 32'd54009;
			11528: outdata = 32'd54008;
			11529: outdata = 32'd54007;
			11530: outdata = 32'd54006;
			11531: outdata = 32'd54005;
			11532: outdata = 32'd54004;
			11533: outdata = 32'd54003;
			11534: outdata = 32'd54002;
			11535: outdata = 32'd54001;
			11536: outdata = 32'd54000;
			11537: outdata = 32'd53999;
			11538: outdata = 32'd53998;
			11539: outdata = 32'd53997;
			11540: outdata = 32'd53996;
			11541: outdata = 32'd53995;
			11542: outdata = 32'd53994;
			11543: outdata = 32'd53993;
			11544: outdata = 32'd53992;
			11545: outdata = 32'd53991;
			11546: outdata = 32'd53990;
			11547: outdata = 32'd53989;
			11548: outdata = 32'd53988;
			11549: outdata = 32'd53987;
			11550: outdata = 32'd53986;
			11551: outdata = 32'd53985;
			11552: outdata = 32'd53984;
			11553: outdata = 32'd53983;
			11554: outdata = 32'd53982;
			11555: outdata = 32'd53981;
			11556: outdata = 32'd53980;
			11557: outdata = 32'd53979;
			11558: outdata = 32'd53978;
			11559: outdata = 32'd53977;
			11560: outdata = 32'd53976;
			11561: outdata = 32'd53975;
			11562: outdata = 32'd53974;
			11563: outdata = 32'd53973;
			11564: outdata = 32'd53972;
			11565: outdata = 32'd53971;
			11566: outdata = 32'd53970;
			11567: outdata = 32'd53969;
			11568: outdata = 32'd53968;
			11569: outdata = 32'd53967;
			11570: outdata = 32'd53966;
			11571: outdata = 32'd53965;
			11572: outdata = 32'd53964;
			11573: outdata = 32'd53963;
			11574: outdata = 32'd53962;
			11575: outdata = 32'd53961;
			11576: outdata = 32'd53960;
			11577: outdata = 32'd53959;
			11578: outdata = 32'd53958;
			11579: outdata = 32'd53957;
			11580: outdata = 32'd53956;
			11581: outdata = 32'd53955;
			11582: outdata = 32'd53954;
			11583: outdata = 32'd53953;
			11584: outdata = 32'd53952;
			11585: outdata = 32'd53951;
			11586: outdata = 32'd53950;
			11587: outdata = 32'd53949;
			11588: outdata = 32'd53948;
			11589: outdata = 32'd53947;
			11590: outdata = 32'd53946;
			11591: outdata = 32'd53945;
			11592: outdata = 32'd53944;
			11593: outdata = 32'd53943;
			11594: outdata = 32'd53942;
			11595: outdata = 32'd53941;
			11596: outdata = 32'd53940;
			11597: outdata = 32'd53939;
			11598: outdata = 32'd53938;
			11599: outdata = 32'd53937;
			11600: outdata = 32'd53936;
			11601: outdata = 32'd53935;
			11602: outdata = 32'd53934;
			11603: outdata = 32'd53933;
			11604: outdata = 32'd53932;
			11605: outdata = 32'd53931;
			11606: outdata = 32'd53930;
			11607: outdata = 32'd53929;
			11608: outdata = 32'd53928;
			11609: outdata = 32'd53927;
			11610: outdata = 32'd53926;
			11611: outdata = 32'd53925;
			11612: outdata = 32'd53924;
			11613: outdata = 32'd53923;
			11614: outdata = 32'd53922;
			11615: outdata = 32'd53921;
			11616: outdata = 32'd53920;
			11617: outdata = 32'd53919;
			11618: outdata = 32'd53918;
			11619: outdata = 32'd53917;
			11620: outdata = 32'd53916;
			11621: outdata = 32'd53915;
			11622: outdata = 32'd53914;
			11623: outdata = 32'd53913;
			11624: outdata = 32'd53912;
			11625: outdata = 32'd53911;
			11626: outdata = 32'd53910;
			11627: outdata = 32'd53909;
			11628: outdata = 32'd53908;
			11629: outdata = 32'd53907;
			11630: outdata = 32'd53906;
			11631: outdata = 32'd53905;
			11632: outdata = 32'd53904;
			11633: outdata = 32'd53903;
			11634: outdata = 32'd53902;
			11635: outdata = 32'd53901;
			11636: outdata = 32'd53900;
			11637: outdata = 32'd53899;
			11638: outdata = 32'd53898;
			11639: outdata = 32'd53897;
			11640: outdata = 32'd53896;
			11641: outdata = 32'd53895;
			11642: outdata = 32'd53894;
			11643: outdata = 32'd53893;
			11644: outdata = 32'd53892;
			11645: outdata = 32'd53891;
			11646: outdata = 32'd53890;
			11647: outdata = 32'd53889;
			11648: outdata = 32'd53888;
			11649: outdata = 32'd53887;
			11650: outdata = 32'd53886;
			11651: outdata = 32'd53885;
			11652: outdata = 32'd53884;
			11653: outdata = 32'd53883;
			11654: outdata = 32'd53882;
			11655: outdata = 32'd53881;
			11656: outdata = 32'd53880;
			11657: outdata = 32'd53879;
			11658: outdata = 32'd53878;
			11659: outdata = 32'd53877;
			11660: outdata = 32'd53876;
			11661: outdata = 32'd53875;
			11662: outdata = 32'd53874;
			11663: outdata = 32'd53873;
			11664: outdata = 32'd53872;
			11665: outdata = 32'd53871;
			11666: outdata = 32'd53870;
			11667: outdata = 32'd53869;
			11668: outdata = 32'd53868;
			11669: outdata = 32'd53867;
			11670: outdata = 32'd53866;
			11671: outdata = 32'd53865;
			11672: outdata = 32'd53864;
			11673: outdata = 32'd53863;
			11674: outdata = 32'd53862;
			11675: outdata = 32'd53861;
			11676: outdata = 32'd53860;
			11677: outdata = 32'd53859;
			11678: outdata = 32'd53858;
			11679: outdata = 32'd53857;
			11680: outdata = 32'd53856;
			11681: outdata = 32'd53855;
			11682: outdata = 32'd53854;
			11683: outdata = 32'd53853;
			11684: outdata = 32'd53852;
			11685: outdata = 32'd53851;
			11686: outdata = 32'd53850;
			11687: outdata = 32'd53849;
			11688: outdata = 32'd53848;
			11689: outdata = 32'd53847;
			11690: outdata = 32'd53846;
			11691: outdata = 32'd53845;
			11692: outdata = 32'd53844;
			11693: outdata = 32'd53843;
			11694: outdata = 32'd53842;
			11695: outdata = 32'd53841;
			11696: outdata = 32'd53840;
			11697: outdata = 32'd53839;
			11698: outdata = 32'd53838;
			11699: outdata = 32'd53837;
			11700: outdata = 32'd53836;
			11701: outdata = 32'd53835;
			11702: outdata = 32'd53834;
			11703: outdata = 32'd53833;
			11704: outdata = 32'd53832;
			11705: outdata = 32'd53831;
			11706: outdata = 32'd53830;
			11707: outdata = 32'd53829;
			11708: outdata = 32'd53828;
			11709: outdata = 32'd53827;
			11710: outdata = 32'd53826;
			11711: outdata = 32'd53825;
			11712: outdata = 32'd53824;
			11713: outdata = 32'd53823;
			11714: outdata = 32'd53822;
			11715: outdata = 32'd53821;
			11716: outdata = 32'd53820;
			11717: outdata = 32'd53819;
			11718: outdata = 32'd53818;
			11719: outdata = 32'd53817;
			11720: outdata = 32'd53816;
			11721: outdata = 32'd53815;
			11722: outdata = 32'd53814;
			11723: outdata = 32'd53813;
			11724: outdata = 32'd53812;
			11725: outdata = 32'd53811;
			11726: outdata = 32'd53810;
			11727: outdata = 32'd53809;
			11728: outdata = 32'd53808;
			11729: outdata = 32'd53807;
			11730: outdata = 32'd53806;
			11731: outdata = 32'd53805;
			11732: outdata = 32'd53804;
			11733: outdata = 32'd53803;
			11734: outdata = 32'd53802;
			11735: outdata = 32'd53801;
			11736: outdata = 32'd53800;
			11737: outdata = 32'd53799;
			11738: outdata = 32'd53798;
			11739: outdata = 32'd53797;
			11740: outdata = 32'd53796;
			11741: outdata = 32'd53795;
			11742: outdata = 32'd53794;
			11743: outdata = 32'd53793;
			11744: outdata = 32'd53792;
			11745: outdata = 32'd53791;
			11746: outdata = 32'd53790;
			11747: outdata = 32'd53789;
			11748: outdata = 32'd53788;
			11749: outdata = 32'd53787;
			11750: outdata = 32'd53786;
			11751: outdata = 32'd53785;
			11752: outdata = 32'd53784;
			11753: outdata = 32'd53783;
			11754: outdata = 32'd53782;
			11755: outdata = 32'd53781;
			11756: outdata = 32'd53780;
			11757: outdata = 32'd53779;
			11758: outdata = 32'd53778;
			11759: outdata = 32'd53777;
			11760: outdata = 32'd53776;
			11761: outdata = 32'd53775;
			11762: outdata = 32'd53774;
			11763: outdata = 32'd53773;
			11764: outdata = 32'd53772;
			11765: outdata = 32'd53771;
			11766: outdata = 32'd53770;
			11767: outdata = 32'd53769;
			11768: outdata = 32'd53768;
			11769: outdata = 32'd53767;
			11770: outdata = 32'd53766;
			11771: outdata = 32'd53765;
			11772: outdata = 32'd53764;
			11773: outdata = 32'd53763;
			11774: outdata = 32'd53762;
			11775: outdata = 32'd53761;
			11776: outdata = 32'd53760;
			11777: outdata = 32'd53759;
			11778: outdata = 32'd53758;
			11779: outdata = 32'd53757;
			11780: outdata = 32'd53756;
			11781: outdata = 32'd53755;
			11782: outdata = 32'd53754;
			11783: outdata = 32'd53753;
			11784: outdata = 32'd53752;
			11785: outdata = 32'd53751;
			11786: outdata = 32'd53750;
			11787: outdata = 32'd53749;
			11788: outdata = 32'd53748;
			11789: outdata = 32'd53747;
			11790: outdata = 32'd53746;
			11791: outdata = 32'd53745;
			11792: outdata = 32'd53744;
			11793: outdata = 32'd53743;
			11794: outdata = 32'd53742;
			11795: outdata = 32'd53741;
			11796: outdata = 32'd53740;
			11797: outdata = 32'd53739;
			11798: outdata = 32'd53738;
			11799: outdata = 32'd53737;
			11800: outdata = 32'd53736;
			11801: outdata = 32'd53735;
			11802: outdata = 32'd53734;
			11803: outdata = 32'd53733;
			11804: outdata = 32'd53732;
			11805: outdata = 32'd53731;
			11806: outdata = 32'd53730;
			11807: outdata = 32'd53729;
			11808: outdata = 32'd53728;
			11809: outdata = 32'd53727;
			11810: outdata = 32'd53726;
			11811: outdata = 32'd53725;
			11812: outdata = 32'd53724;
			11813: outdata = 32'd53723;
			11814: outdata = 32'd53722;
			11815: outdata = 32'd53721;
			11816: outdata = 32'd53720;
			11817: outdata = 32'd53719;
			11818: outdata = 32'd53718;
			11819: outdata = 32'd53717;
			11820: outdata = 32'd53716;
			11821: outdata = 32'd53715;
			11822: outdata = 32'd53714;
			11823: outdata = 32'd53713;
			11824: outdata = 32'd53712;
			11825: outdata = 32'd53711;
			11826: outdata = 32'd53710;
			11827: outdata = 32'd53709;
			11828: outdata = 32'd53708;
			11829: outdata = 32'd53707;
			11830: outdata = 32'd53706;
			11831: outdata = 32'd53705;
			11832: outdata = 32'd53704;
			11833: outdata = 32'd53703;
			11834: outdata = 32'd53702;
			11835: outdata = 32'd53701;
			11836: outdata = 32'd53700;
			11837: outdata = 32'd53699;
			11838: outdata = 32'd53698;
			11839: outdata = 32'd53697;
			11840: outdata = 32'd53696;
			11841: outdata = 32'd53695;
			11842: outdata = 32'd53694;
			11843: outdata = 32'd53693;
			11844: outdata = 32'd53692;
			11845: outdata = 32'd53691;
			11846: outdata = 32'd53690;
			11847: outdata = 32'd53689;
			11848: outdata = 32'd53688;
			11849: outdata = 32'd53687;
			11850: outdata = 32'd53686;
			11851: outdata = 32'd53685;
			11852: outdata = 32'd53684;
			11853: outdata = 32'd53683;
			11854: outdata = 32'd53682;
			11855: outdata = 32'd53681;
			11856: outdata = 32'd53680;
			11857: outdata = 32'd53679;
			11858: outdata = 32'd53678;
			11859: outdata = 32'd53677;
			11860: outdata = 32'd53676;
			11861: outdata = 32'd53675;
			11862: outdata = 32'd53674;
			11863: outdata = 32'd53673;
			11864: outdata = 32'd53672;
			11865: outdata = 32'd53671;
			11866: outdata = 32'd53670;
			11867: outdata = 32'd53669;
			11868: outdata = 32'd53668;
			11869: outdata = 32'd53667;
			11870: outdata = 32'd53666;
			11871: outdata = 32'd53665;
			11872: outdata = 32'd53664;
			11873: outdata = 32'd53663;
			11874: outdata = 32'd53662;
			11875: outdata = 32'd53661;
			11876: outdata = 32'd53660;
			11877: outdata = 32'd53659;
			11878: outdata = 32'd53658;
			11879: outdata = 32'd53657;
			11880: outdata = 32'd53656;
			11881: outdata = 32'd53655;
			11882: outdata = 32'd53654;
			11883: outdata = 32'd53653;
			11884: outdata = 32'd53652;
			11885: outdata = 32'd53651;
			11886: outdata = 32'd53650;
			11887: outdata = 32'd53649;
			11888: outdata = 32'd53648;
			11889: outdata = 32'd53647;
			11890: outdata = 32'd53646;
			11891: outdata = 32'd53645;
			11892: outdata = 32'd53644;
			11893: outdata = 32'd53643;
			11894: outdata = 32'd53642;
			11895: outdata = 32'd53641;
			11896: outdata = 32'd53640;
			11897: outdata = 32'd53639;
			11898: outdata = 32'd53638;
			11899: outdata = 32'd53637;
			11900: outdata = 32'd53636;
			11901: outdata = 32'd53635;
			11902: outdata = 32'd53634;
			11903: outdata = 32'd53633;
			11904: outdata = 32'd53632;
			11905: outdata = 32'd53631;
			11906: outdata = 32'd53630;
			11907: outdata = 32'd53629;
			11908: outdata = 32'd53628;
			11909: outdata = 32'd53627;
			11910: outdata = 32'd53626;
			11911: outdata = 32'd53625;
			11912: outdata = 32'd53624;
			11913: outdata = 32'd53623;
			11914: outdata = 32'd53622;
			11915: outdata = 32'd53621;
			11916: outdata = 32'd53620;
			11917: outdata = 32'd53619;
			11918: outdata = 32'd53618;
			11919: outdata = 32'd53617;
			11920: outdata = 32'd53616;
			11921: outdata = 32'd53615;
			11922: outdata = 32'd53614;
			11923: outdata = 32'd53613;
			11924: outdata = 32'd53612;
			11925: outdata = 32'd53611;
			11926: outdata = 32'd53610;
			11927: outdata = 32'd53609;
			11928: outdata = 32'd53608;
			11929: outdata = 32'd53607;
			11930: outdata = 32'd53606;
			11931: outdata = 32'd53605;
			11932: outdata = 32'd53604;
			11933: outdata = 32'd53603;
			11934: outdata = 32'd53602;
			11935: outdata = 32'd53601;
			11936: outdata = 32'd53600;
			11937: outdata = 32'd53599;
			11938: outdata = 32'd53598;
			11939: outdata = 32'd53597;
			11940: outdata = 32'd53596;
			11941: outdata = 32'd53595;
			11942: outdata = 32'd53594;
			11943: outdata = 32'd53593;
			11944: outdata = 32'd53592;
			11945: outdata = 32'd53591;
			11946: outdata = 32'd53590;
			11947: outdata = 32'd53589;
			11948: outdata = 32'd53588;
			11949: outdata = 32'd53587;
			11950: outdata = 32'd53586;
			11951: outdata = 32'd53585;
			11952: outdata = 32'd53584;
			11953: outdata = 32'd53583;
			11954: outdata = 32'd53582;
			11955: outdata = 32'd53581;
			11956: outdata = 32'd53580;
			11957: outdata = 32'd53579;
			11958: outdata = 32'd53578;
			11959: outdata = 32'd53577;
			11960: outdata = 32'd53576;
			11961: outdata = 32'd53575;
			11962: outdata = 32'd53574;
			11963: outdata = 32'd53573;
			11964: outdata = 32'd53572;
			11965: outdata = 32'd53571;
			11966: outdata = 32'd53570;
			11967: outdata = 32'd53569;
			11968: outdata = 32'd53568;
			11969: outdata = 32'd53567;
			11970: outdata = 32'd53566;
			11971: outdata = 32'd53565;
			11972: outdata = 32'd53564;
			11973: outdata = 32'd53563;
			11974: outdata = 32'd53562;
			11975: outdata = 32'd53561;
			11976: outdata = 32'd53560;
			11977: outdata = 32'd53559;
			11978: outdata = 32'd53558;
			11979: outdata = 32'd53557;
			11980: outdata = 32'd53556;
			11981: outdata = 32'd53555;
			11982: outdata = 32'd53554;
			11983: outdata = 32'd53553;
			11984: outdata = 32'd53552;
			11985: outdata = 32'd53551;
			11986: outdata = 32'd53550;
			11987: outdata = 32'd53549;
			11988: outdata = 32'd53548;
			11989: outdata = 32'd53547;
			11990: outdata = 32'd53546;
			11991: outdata = 32'd53545;
			11992: outdata = 32'd53544;
			11993: outdata = 32'd53543;
			11994: outdata = 32'd53542;
			11995: outdata = 32'd53541;
			11996: outdata = 32'd53540;
			11997: outdata = 32'd53539;
			11998: outdata = 32'd53538;
			11999: outdata = 32'd53537;
			12000: outdata = 32'd53536;
			12001: outdata = 32'd53535;
			12002: outdata = 32'd53534;
			12003: outdata = 32'd53533;
			12004: outdata = 32'd53532;
			12005: outdata = 32'd53531;
			12006: outdata = 32'd53530;
			12007: outdata = 32'd53529;
			12008: outdata = 32'd53528;
			12009: outdata = 32'd53527;
			12010: outdata = 32'd53526;
			12011: outdata = 32'd53525;
			12012: outdata = 32'd53524;
			12013: outdata = 32'd53523;
			12014: outdata = 32'd53522;
			12015: outdata = 32'd53521;
			12016: outdata = 32'd53520;
			12017: outdata = 32'd53519;
			12018: outdata = 32'd53518;
			12019: outdata = 32'd53517;
			12020: outdata = 32'd53516;
			12021: outdata = 32'd53515;
			12022: outdata = 32'd53514;
			12023: outdata = 32'd53513;
			12024: outdata = 32'd53512;
			12025: outdata = 32'd53511;
			12026: outdata = 32'd53510;
			12027: outdata = 32'd53509;
			12028: outdata = 32'd53508;
			12029: outdata = 32'd53507;
			12030: outdata = 32'd53506;
			12031: outdata = 32'd53505;
			12032: outdata = 32'd53504;
			12033: outdata = 32'd53503;
			12034: outdata = 32'd53502;
			12035: outdata = 32'd53501;
			12036: outdata = 32'd53500;
			12037: outdata = 32'd53499;
			12038: outdata = 32'd53498;
			12039: outdata = 32'd53497;
			12040: outdata = 32'd53496;
			12041: outdata = 32'd53495;
			12042: outdata = 32'd53494;
			12043: outdata = 32'd53493;
			12044: outdata = 32'd53492;
			12045: outdata = 32'd53491;
			12046: outdata = 32'd53490;
			12047: outdata = 32'd53489;
			12048: outdata = 32'd53488;
			12049: outdata = 32'd53487;
			12050: outdata = 32'd53486;
			12051: outdata = 32'd53485;
			12052: outdata = 32'd53484;
			12053: outdata = 32'd53483;
			12054: outdata = 32'd53482;
			12055: outdata = 32'd53481;
			12056: outdata = 32'd53480;
			12057: outdata = 32'd53479;
			12058: outdata = 32'd53478;
			12059: outdata = 32'd53477;
			12060: outdata = 32'd53476;
			12061: outdata = 32'd53475;
			12062: outdata = 32'd53474;
			12063: outdata = 32'd53473;
			12064: outdata = 32'd53472;
			12065: outdata = 32'd53471;
			12066: outdata = 32'd53470;
			12067: outdata = 32'd53469;
			12068: outdata = 32'd53468;
			12069: outdata = 32'd53467;
			12070: outdata = 32'd53466;
			12071: outdata = 32'd53465;
			12072: outdata = 32'd53464;
			12073: outdata = 32'd53463;
			12074: outdata = 32'd53462;
			12075: outdata = 32'd53461;
			12076: outdata = 32'd53460;
			12077: outdata = 32'd53459;
			12078: outdata = 32'd53458;
			12079: outdata = 32'd53457;
			12080: outdata = 32'd53456;
			12081: outdata = 32'd53455;
			12082: outdata = 32'd53454;
			12083: outdata = 32'd53453;
			12084: outdata = 32'd53452;
			12085: outdata = 32'd53451;
			12086: outdata = 32'd53450;
			12087: outdata = 32'd53449;
			12088: outdata = 32'd53448;
			12089: outdata = 32'd53447;
			12090: outdata = 32'd53446;
			12091: outdata = 32'd53445;
			12092: outdata = 32'd53444;
			12093: outdata = 32'd53443;
			12094: outdata = 32'd53442;
			12095: outdata = 32'd53441;
			12096: outdata = 32'd53440;
			12097: outdata = 32'd53439;
			12098: outdata = 32'd53438;
			12099: outdata = 32'd53437;
			12100: outdata = 32'd53436;
			12101: outdata = 32'd53435;
			12102: outdata = 32'd53434;
			12103: outdata = 32'd53433;
			12104: outdata = 32'd53432;
			12105: outdata = 32'd53431;
			12106: outdata = 32'd53430;
			12107: outdata = 32'd53429;
			12108: outdata = 32'd53428;
			12109: outdata = 32'd53427;
			12110: outdata = 32'd53426;
			12111: outdata = 32'd53425;
			12112: outdata = 32'd53424;
			12113: outdata = 32'd53423;
			12114: outdata = 32'd53422;
			12115: outdata = 32'd53421;
			12116: outdata = 32'd53420;
			12117: outdata = 32'd53419;
			12118: outdata = 32'd53418;
			12119: outdata = 32'd53417;
			12120: outdata = 32'd53416;
			12121: outdata = 32'd53415;
			12122: outdata = 32'd53414;
			12123: outdata = 32'd53413;
			12124: outdata = 32'd53412;
			12125: outdata = 32'd53411;
			12126: outdata = 32'd53410;
			12127: outdata = 32'd53409;
			12128: outdata = 32'd53408;
			12129: outdata = 32'd53407;
			12130: outdata = 32'd53406;
			12131: outdata = 32'd53405;
			12132: outdata = 32'd53404;
			12133: outdata = 32'd53403;
			12134: outdata = 32'd53402;
			12135: outdata = 32'd53401;
			12136: outdata = 32'd53400;
			12137: outdata = 32'd53399;
			12138: outdata = 32'd53398;
			12139: outdata = 32'd53397;
			12140: outdata = 32'd53396;
			12141: outdata = 32'd53395;
			12142: outdata = 32'd53394;
			12143: outdata = 32'd53393;
			12144: outdata = 32'd53392;
			12145: outdata = 32'd53391;
			12146: outdata = 32'd53390;
			12147: outdata = 32'd53389;
			12148: outdata = 32'd53388;
			12149: outdata = 32'd53387;
			12150: outdata = 32'd53386;
			12151: outdata = 32'd53385;
			12152: outdata = 32'd53384;
			12153: outdata = 32'd53383;
			12154: outdata = 32'd53382;
			12155: outdata = 32'd53381;
			12156: outdata = 32'd53380;
			12157: outdata = 32'd53379;
			12158: outdata = 32'd53378;
			12159: outdata = 32'd53377;
			12160: outdata = 32'd53376;
			12161: outdata = 32'd53375;
			12162: outdata = 32'd53374;
			12163: outdata = 32'd53373;
			12164: outdata = 32'd53372;
			12165: outdata = 32'd53371;
			12166: outdata = 32'd53370;
			12167: outdata = 32'd53369;
			12168: outdata = 32'd53368;
			12169: outdata = 32'd53367;
			12170: outdata = 32'd53366;
			12171: outdata = 32'd53365;
			12172: outdata = 32'd53364;
			12173: outdata = 32'd53363;
			12174: outdata = 32'd53362;
			12175: outdata = 32'd53361;
			12176: outdata = 32'd53360;
			12177: outdata = 32'd53359;
			12178: outdata = 32'd53358;
			12179: outdata = 32'd53357;
			12180: outdata = 32'd53356;
			12181: outdata = 32'd53355;
			12182: outdata = 32'd53354;
			12183: outdata = 32'd53353;
			12184: outdata = 32'd53352;
			12185: outdata = 32'd53351;
			12186: outdata = 32'd53350;
			12187: outdata = 32'd53349;
			12188: outdata = 32'd53348;
			12189: outdata = 32'd53347;
			12190: outdata = 32'd53346;
			12191: outdata = 32'd53345;
			12192: outdata = 32'd53344;
			12193: outdata = 32'd53343;
			12194: outdata = 32'd53342;
			12195: outdata = 32'd53341;
			12196: outdata = 32'd53340;
			12197: outdata = 32'd53339;
			12198: outdata = 32'd53338;
			12199: outdata = 32'd53337;
			12200: outdata = 32'd53336;
			12201: outdata = 32'd53335;
			12202: outdata = 32'd53334;
			12203: outdata = 32'd53333;
			12204: outdata = 32'd53332;
			12205: outdata = 32'd53331;
			12206: outdata = 32'd53330;
			12207: outdata = 32'd53329;
			12208: outdata = 32'd53328;
			12209: outdata = 32'd53327;
			12210: outdata = 32'd53326;
			12211: outdata = 32'd53325;
			12212: outdata = 32'd53324;
			12213: outdata = 32'd53323;
			12214: outdata = 32'd53322;
			12215: outdata = 32'd53321;
			12216: outdata = 32'd53320;
			12217: outdata = 32'd53319;
			12218: outdata = 32'd53318;
			12219: outdata = 32'd53317;
			12220: outdata = 32'd53316;
			12221: outdata = 32'd53315;
			12222: outdata = 32'd53314;
			12223: outdata = 32'd53313;
			12224: outdata = 32'd53312;
			12225: outdata = 32'd53311;
			12226: outdata = 32'd53310;
			12227: outdata = 32'd53309;
			12228: outdata = 32'd53308;
			12229: outdata = 32'd53307;
			12230: outdata = 32'd53306;
			12231: outdata = 32'd53305;
			12232: outdata = 32'd53304;
			12233: outdata = 32'd53303;
			12234: outdata = 32'd53302;
			12235: outdata = 32'd53301;
			12236: outdata = 32'd53300;
			12237: outdata = 32'd53299;
			12238: outdata = 32'd53298;
			12239: outdata = 32'd53297;
			12240: outdata = 32'd53296;
			12241: outdata = 32'd53295;
			12242: outdata = 32'd53294;
			12243: outdata = 32'd53293;
			12244: outdata = 32'd53292;
			12245: outdata = 32'd53291;
			12246: outdata = 32'd53290;
			12247: outdata = 32'd53289;
			12248: outdata = 32'd53288;
			12249: outdata = 32'd53287;
			12250: outdata = 32'd53286;
			12251: outdata = 32'd53285;
			12252: outdata = 32'd53284;
			12253: outdata = 32'd53283;
			12254: outdata = 32'd53282;
			12255: outdata = 32'd53281;
			12256: outdata = 32'd53280;
			12257: outdata = 32'd53279;
			12258: outdata = 32'd53278;
			12259: outdata = 32'd53277;
			12260: outdata = 32'd53276;
			12261: outdata = 32'd53275;
			12262: outdata = 32'd53274;
			12263: outdata = 32'd53273;
			12264: outdata = 32'd53272;
			12265: outdata = 32'd53271;
			12266: outdata = 32'd53270;
			12267: outdata = 32'd53269;
			12268: outdata = 32'd53268;
			12269: outdata = 32'd53267;
			12270: outdata = 32'd53266;
			12271: outdata = 32'd53265;
			12272: outdata = 32'd53264;
			12273: outdata = 32'd53263;
			12274: outdata = 32'd53262;
			12275: outdata = 32'd53261;
			12276: outdata = 32'd53260;
			12277: outdata = 32'd53259;
			12278: outdata = 32'd53258;
			12279: outdata = 32'd53257;
			12280: outdata = 32'd53256;
			12281: outdata = 32'd53255;
			12282: outdata = 32'd53254;
			12283: outdata = 32'd53253;
			12284: outdata = 32'd53252;
			12285: outdata = 32'd53251;
			12286: outdata = 32'd53250;
			12287: outdata = 32'd53249;
			12288: outdata = 32'd53248;
			12289: outdata = 32'd53247;
			12290: outdata = 32'd53246;
			12291: outdata = 32'd53245;
			12292: outdata = 32'd53244;
			12293: outdata = 32'd53243;
			12294: outdata = 32'd53242;
			12295: outdata = 32'd53241;
			12296: outdata = 32'd53240;
			12297: outdata = 32'd53239;
			12298: outdata = 32'd53238;
			12299: outdata = 32'd53237;
			12300: outdata = 32'd53236;
			12301: outdata = 32'd53235;
			12302: outdata = 32'd53234;
			12303: outdata = 32'd53233;
			12304: outdata = 32'd53232;
			12305: outdata = 32'd53231;
			12306: outdata = 32'd53230;
			12307: outdata = 32'd53229;
			12308: outdata = 32'd53228;
			12309: outdata = 32'd53227;
			12310: outdata = 32'd53226;
			12311: outdata = 32'd53225;
			12312: outdata = 32'd53224;
			12313: outdata = 32'd53223;
			12314: outdata = 32'd53222;
			12315: outdata = 32'd53221;
			12316: outdata = 32'd53220;
			12317: outdata = 32'd53219;
			12318: outdata = 32'd53218;
			12319: outdata = 32'd53217;
			12320: outdata = 32'd53216;
			12321: outdata = 32'd53215;
			12322: outdata = 32'd53214;
			12323: outdata = 32'd53213;
			12324: outdata = 32'd53212;
			12325: outdata = 32'd53211;
			12326: outdata = 32'd53210;
			12327: outdata = 32'd53209;
			12328: outdata = 32'd53208;
			12329: outdata = 32'd53207;
			12330: outdata = 32'd53206;
			12331: outdata = 32'd53205;
			12332: outdata = 32'd53204;
			12333: outdata = 32'd53203;
			12334: outdata = 32'd53202;
			12335: outdata = 32'd53201;
			12336: outdata = 32'd53200;
			12337: outdata = 32'd53199;
			12338: outdata = 32'd53198;
			12339: outdata = 32'd53197;
			12340: outdata = 32'd53196;
			12341: outdata = 32'd53195;
			12342: outdata = 32'd53194;
			12343: outdata = 32'd53193;
			12344: outdata = 32'd53192;
			12345: outdata = 32'd53191;
			12346: outdata = 32'd53190;
			12347: outdata = 32'd53189;
			12348: outdata = 32'd53188;
			12349: outdata = 32'd53187;
			12350: outdata = 32'd53186;
			12351: outdata = 32'd53185;
			12352: outdata = 32'd53184;
			12353: outdata = 32'd53183;
			12354: outdata = 32'd53182;
			12355: outdata = 32'd53181;
			12356: outdata = 32'd53180;
			12357: outdata = 32'd53179;
			12358: outdata = 32'd53178;
			12359: outdata = 32'd53177;
			12360: outdata = 32'd53176;
			12361: outdata = 32'd53175;
			12362: outdata = 32'd53174;
			12363: outdata = 32'd53173;
			12364: outdata = 32'd53172;
			12365: outdata = 32'd53171;
			12366: outdata = 32'd53170;
			12367: outdata = 32'd53169;
			12368: outdata = 32'd53168;
			12369: outdata = 32'd53167;
			12370: outdata = 32'd53166;
			12371: outdata = 32'd53165;
			12372: outdata = 32'd53164;
			12373: outdata = 32'd53163;
			12374: outdata = 32'd53162;
			12375: outdata = 32'd53161;
			12376: outdata = 32'd53160;
			12377: outdata = 32'd53159;
			12378: outdata = 32'd53158;
			12379: outdata = 32'd53157;
			12380: outdata = 32'd53156;
			12381: outdata = 32'd53155;
			12382: outdata = 32'd53154;
			12383: outdata = 32'd53153;
			12384: outdata = 32'd53152;
			12385: outdata = 32'd53151;
			12386: outdata = 32'd53150;
			12387: outdata = 32'd53149;
			12388: outdata = 32'd53148;
			12389: outdata = 32'd53147;
			12390: outdata = 32'd53146;
			12391: outdata = 32'd53145;
			12392: outdata = 32'd53144;
			12393: outdata = 32'd53143;
			12394: outdata = 32'd53142;
			12395: outdata = 32'd53141;
			12396: outdata = 32'd53140;
			12397: outdata = 32'd53139;
			12398: outdata = 32'd53138;
			12399: outdata = 32'd53137;
			12400: outdata = 32'd53136;
			12401: outdata = 32'd53135;
			12402: outdata = 32'd53134;
			12403: outdata = 32'd53133;
			12404: outdata = 32'd53132;
			12405: outdata = 32'd53131;
			12406: outdata = 32'd53130;
			12407: outdata = 32'd53129;
			12408: outdata = 32'd53128;
			12409: outdata = 32'd53127;
			12410: outdata = 32'd53126;
			12411: outdata = 32'd53125;
			12412: outdata = 32'd53124;
			12413: outdata = 32'd53123;
			12414: outdata = 32'd53122;
			12415: outdata = 32'd53121;
			12416: outdata = 32'd53120;
			12417: outdata = 32'd53119;
			12418: outdata = 32'd53118;
			12419: outdata = 32'd53117;
			12420: outdata = 32'd53116;
			12421: outdata = 32'd53115;
			12422: outdata = 32'd53114;
			12423: outdata = 32'd53113;
			12424: outdata = 32'd53112;
			12425: outdata = 32'd53111;
			12426: outdata = 32'd53110;
			12427: outdata = 32'd53109;
			12428: outdata = 32'd53108;
			12429: outdata = 32'd53107;
			12430: outdata = 32'd53106;
			12431: outdata = 32'd53105;
			12432: outdata = 32'd53104;
			12433: outdata = 32'd53103;
			12434: outdata = 32'd53102;
			12435: outdata = 32'd53101;
			12436: outdata = 32'd53100;
			12437: outdata = 32'd53099;
			12438: outdata = 32'd53098;
			12439: outdata = 32'd53097;
			12440: outdata = 32'd53096;
			12441: outdata = 32'd53095;
			12442: outdata = 32'd53094;
			12443: outdata = 32'd53093;
			12444: outdata = 32'd53092;
			12445: outdata = 32'd53091;
			12446: outdata = 32'd53090;
			12447: outdata = 32'd53089;
			12448: outdata = 32'd53088;
			12449: outdata = 32'd53087;
			12450: outdata = 32'd53086;
			12451: outdata = 32'd53085;
			12452: outdata = 32'd53084;
			12453: outdata = 32'd53083;
			12454: outdata = 32'd53082;
			12455: outdata = 32'd53081;
			12456: outdata = 32'd53080;
			12457: outdata = 32'd53079;
			12458: outdata = 32'd53078;
			12459: outdata = 32'd53077;
			12460: outdata = 32'd53076;
			12461: outdata = 32'd53075;
			12462: outdata = 32'd53074;
			12463: outdata = 32'd53073;
			12464: outdata = 32'd53072;
			12465: outdata = 32'd53071;
			12466: outdata = 32'd53070;
			12467: outdata = 32'd53069;
			12468: outdata = 32'd53068;
			12469: outdata = 32'd53067;
			12470: outdata = 32'd53066;
			12471: outdata = 32'd53065;
			12472: outdata = 32'd53064;
			12473: outdata = 32'd53063;
			12474: outdata = 32'd53062;
			12475: outdata = 32'd53061;
			12476: outdata = 32'd53060;
			12477: outdata = 32'd53059;
			12478: outdata = 32'd53058;
			12479: outdata = 32'd53057;
			12480: outdata = 32'd53056;
			12481: outdata = 32'd53055;
			12482: outdata = 32'd53054;
			12483: outdata = 32'd53053;
			12484: outdata = 32'd53052;
			12485: outdata = 32'd53051;
			12486: outdata = 32'd53050;
			12487: outdata = 32'd53049;
			12488: outdata = 32'd53048;
			12489: outdata = 32'd53047;
			12490: outdata = 32'd53046;
			12491: outdata = 32'd53045;
			12492: outdata = 32'd53044;
			12493: outdata = 32'd53043;
			12494: outdata = 32'd53042;
			12495: outdata = 32'd53041;
			12496: outdata = 32'd53040;
			12497: outdata = 32'd53039;
			12498: outdata = 32'd53038;
			12499: outdata = 32'd53037;
			12500: outdata = 32'd53036;
			12501: outdata = 32'd53035;
			12502: outdata = 32'd53034;
			12503: outdata = 32'd53033;
			12504: outdata = 32'd53032;
			12505: outdata = 32'd53031;
			12506: outdata = 32'd53030;
			12507: outdata = 32'd53029;
			12508: outdata = 32'd53028;
			12509: outdata = 32'd53027;
			12510: outdata = 32'd53026;
			12511: outdata = 32'd53025;
			12512: outdata = 32'd53024;
			12513: outdata = 32'd53023;
			12514: outdata = 32'd53022;
			12515: outdata = 32'd53021;
			12516: outdata = 32'd53020;
			12517: outdata = 32'd53019;
			12518: outdata = 32'd53018;
			12519: outdata = 32'd53017;
			12520: outdata = 32'd53016;
			12521: outdata = 32'd53015;
			12522: outdata = 32'd53014;
			12523: outdata = 32'd53013;
			12524: outdata = 32'd53012;
			12525: outdata = 32'd53011;
			12526: outdata = 32'd53010;
			12527: outdata = 32'd53009;
			12528: outdata = 32'd53008;
			12529: outdata = 32'd53007;
			12530: outdata = 32'd53006;
			12531: outdata = 32'd53005;
			12532: outdata = 32'd53004;
			12533: outdata = 32'd53003;
			12534: outdata = 32'd53002;
			12535: outdata = 32'd53001;
			12536: outdata = 32'd53000;
			12537: outdata = 32'd52999;
			12538: outdata = 32'd52998;
			12539: outdata = 32'd52997;
			12540: outdata = 32'd52996;
			12541: outdata = 32'd52995;
			12542: outdata = 32'd52994;
			12543: outdata = 32'd52993;
			12544: outdata = 32'd52992;
			12545: outdata = 32'd52991;
			12546: outdata = 32'd52990;
			12547: outdata = 32'd52989;
			12548: outdata = 32'd52988;
			12549: outdata = 32'd52987;
			12550: outdata = 32'd52986;
			12551: outdata = 32'd52985;
			12552: outdata = 32'd52984;
			12553: outdata = 32'd52983;
			12554: outdata = 32'd52982;
			12555: outdata = 32'd52981;
			12556: outdata = 32'd52980;
			12557: outdata = 32'd52979;
			12558: outdata = 32'd52978;
			12559: outdata = 32'd52977;
			12560: outdata = 32'd52976;
			12561: outdata = 32'd52975;
			12562: outdata = 32'd52974;
			12563: outdata = 32'd52973;
			12564: outdata = 32'd52972;
			12565: outdata = 32'd52971;
			12566: outdata = 32'd52970;
			12567: outdata = 32'd52969;
			12568: outdata = 32'd52968;
			12569: outdata = 32'd52967;
			12570: outdata = 32'd52966;
			12571: outdata = 32'd52965;
			12572: outdata = 32'd52964;
			12573: outdata = 32'd52963;
			12574: outdata = 32'd52962;
			12575: outdata = 32'd52961;
			12576: outdata = 32'd52960;
			12577: outdata = 32'd52959;
			12578: outdata = 32'd52958;
			12579: outdata = 32'd52957;
			12580: outdata = 32'd52956;
			12581: outdata = 32'd52955;
			12582: outdata = 32'd52954;
			12583: outdata = 32'd52953;
			12584: outdata = 32'd52952;
			12585: outdata = 32'd52951;
			12586: outdata = 32'd52950;
			12587: outdata = 32'd52949;
			12588: outdata = 32'd52948;
			12589: outdata = 32'd52947;
			12590: outdata = 32'd52946;
			12591: outdata = 32'd52945;
			12592: outdata = 32'd52944;
			12593: outdata = 32'd52943;
			12594: outdata = 32'd52942;
			12595: outdata = 32'd52941;
			12596: outdata = 32'd52940;
			12597: outdata = 32'd52939;
			12598: outdata = 32'd52938;
			12599: outdata = 32'd52937;
			12600: outdata = 32'd52936;
			12601: outdata = 32'd52935;
			12602: outdata = 32'd52934;
			12603: outdata = 32'd52933;
			12604: outdata = 32'd52932;
			12605: outdata = 32'd52931;
			12606: outdata = 32'd52930;
			12607: outdata = 32'd52929;
			12608: outdata = 32'd52928;
			12609: outdata = 32'd52927;
			12610: outdata = 32'd52926;
			12611: outdata = 32'd52925;
			12612: outdata = 32'd52924;
			12613: outdata = 32'd52923;
			12614: outdata = 32'd52922;
			12615: outdata = 32'd52921;
			12616: outdata = 32'd52920;
			12617: outdata = 32'd52919;
			12618: outdata = 32'd52918;
			12619: outdata = 32'd52917;
			12620: outdata = 32'd52916;
			12621: outdata = 32'd52915;
			12622: outdata = 32'd52914;
			12623: outdata = 32'd52913;
			12624: outdata = 32'd52912;
			12625: outdata = 32'd52911;
			12626: outdata = 32'd52910;
			12627: outdata = 32'd52909;
			12628: outdata = 32'd52908;
			12629: outdata = 32'd52907;
			12630: outdata = 32'd52906;
			12631: outdata = 32'd52905;
			12632: outdata = 32'd52904;
			12633: outdata = 32'd52903;
			12634: outdata = 32'd52902;
			12635: outdata = 32'd52901;
			12636: outdata = 32'd52900;
			12637: outdata = 32'd52899;
			12638: outdata = 32'd52898;
			12639: outdata = 32'd52897;
			12640: outdata = 32'd52896;
			12641: outdata = 32'd52895;
			12642: outdata = 32'd52894;
			12643: outdata = 32'd52893;
			12644: outdata = 32'd52892;
			12645: outdata = 32'd52891;
			12646: outdata = 32'd52890;
			12647: outdata = 32'd52889;
			12648: outdata = 32'd52888;
			12649: outdata = 32'd52887;
			12650: outdata = 32'd52886;
			12651: outdata = 32'd52885;
			12652: outdata = 32'd52884;
			12653: outdata = 32'd52883;
			12654: outdata = 32'd52882;
			12655: outdata = 32'd52881;
			12656: outdata = 32'd52880;
			12657: outdata = 32'd52879;
			12658: outdata = 32'd52878;
			12659: outdata = 32'd52877;
			12660: outdata = 32'd52876;
			12661: outdata = 32'd52875;
			12662: outdata = 32'd52874;
			12663: outdata = 32'd52873;
			12664: outdata = 32'd52872;
			12665: outdata = 32'd52871;
			12666: outdata = 32'd52870;
			12667: outdata = 32'd52869;
			12668: outdata = 32'd52868;
			12669: outdata = 32'd52867;
			12670: outdata = 32'd52866;
			12671: outdata = 32'd52865;
			12672: outdata = 32'd52864;
			12673: outdata = 32'd52863;
			12674: outdata = 32'd52862;
			12675: outdata = 32'd52861;
			12676: outdata = 32'd52860;
			12677: outdata = 32'd52859;
			12678: outdata = 32'd52858;
			12679: outdata = 32'd52857;
			12680: outdata = 32'd52856;
			12681: outdata = 32'd52855;
			12682: outdata = 32'd52854;
			12683: outdata = 32'd52853;
			12684: outdata = 32'd52852;
			12685: outdata = 32'd52851;
			12686: outdata = 32'd52850;
			12687: outdata = 32'd52849;
			12688: outdata = 32'd52848;
			12689: outdata = 32'd52847;
			12690: outdata = 32'd52846;
			12691: outdata = 32'd52845;
			12692: outdata = 32'd52844;
			12693: outdata = 32'd52843;
			12694: outdata = 32'd52842;
			12695: outdata = 32'd52841;
			12696: outdata = 32'd52840;
			12697: outdata = 32'd52839;
			12698: outdata = 32'd52838;
			12699: outdata = 32'd52837;
			12700: outdata = 32'd52836;
			12701: outdata = 32'd52835;
			12702: outdata = 32'd52834;
			12703: outdata = 32'd52833;
			12704: outdata = 32'd52832;
			12705: outdata = 32'd52831;
			12706: outdata = 32'd52830;
			12707: outdata = 32'd52829;
			12708: outdata = 32'd52828;
			12709: outdata = 32'd52827;
			12710: outdata = 32'd52826;
			12711: outdata = 32'd52825;
			12712: outdata = 32'd52824;
			12713: outdata = 32'd52823;
			12714: outdata = 32'd52822;
			12715: outdata = 32'd52821;
			12716: outdata = 32'd52820;
			12717: outdata = 32'd52819;
			12718: outdata = 32'd52818;
			12719: outdata = 32'd52817;
			12720: outdata = 32'd52816;
			12721: outdata = 32'd52815;
			12722: outdata = 32'd52814;
			12723: outdata = 32'd52813;
			12724: outdata = 32'd52812;
			12725: outdata = 32'd52811;
			12726: outdata = 32'd52810;
			12727: outdata = 32'd52809;
			12728: outdata = 32'd52808;
			12729: outdata = 32'd52807;
			12730: outdata = 32'd52806;
			12731: outdata = 32'd52805;
			12732: outdata = 32'd52804;
			12733: outdata = 32'd52803;
			12734: outdata = 32'd52802;
			12735: outdata = 32'd52801;
			12736: outdata = 32'd52800;
			12737: outdata = 32'd52799;
			12738: outdata = 32'd52798;
			12739: outdata = 32'd52797;
			12740: outdata = 32'd52796;
			12741: outdata = 32'd52795;
			12742: outdata = 32'd52794;
			12743: outdata = 32'd52793;
			12744: outdata = 32'd52792;
			12745: outdata = 32'd52791;
			12746: outdata = 32'd52790;
			12747: outdata = 32'd52789;
			12748: outdata = 32'd52788;
			12749: outdata = 32'd52787;
			12750: outdata = 32'd52786;
			12751: outdata = 32'd52785;
			12752: outdata = 32'd52784;
			12753: outdata = 32'd52783;
			12754: outdata = 32'd52782;
			12755: outdata = 32'd52781;
			12756: outdata = 32'd52780;
			12757: outdata = 32'd52779;
			12758: outdata = 32'd52778;
			12759: outdata = 32'd52777;
			12760: outdata = 32'd52776;
			12761: outdata = 32'd52775;
			12762: outdata = 32'd52774;
			12763: outdata = 32'd52773;
			12764: outdata = 32'd52772;
			12765: outdata = 32'd52771;
			12766: outdata = 32'd52770;
			12767: outdata = 32'd52769;
			12768: outdata = 32'd52768;
			12769: outdata = 32'd52767;
			12770: outdata = 32'd52766;
			12771: outdata = 32'd52765;
			12772: outdata = 32'd52764;
			12773: outdata = 32'd52763;
			12774: outdata = 32'd52762;
			12775: outdata = 32'd52761;
			12776: outdata = 32'd52760;
			12777: outdata = 32'd52759;
			12778: outdata = 32'd52758;
			12779: outdata = 32'd52757;
			12780: outdata = 32'd52756;
			12781: outdata = 32'd52755;
			12782: outdata = 32'd52754;
			12783: outdata = 32'd52753;
			12784: outdata = 32'd52752;
			12785: outdata = 32'd52751;
			12786: outdata = 32'd52750;
			12787: outdata = 32'd52749;
			12788: outdata = 32'd52748;
			12789: outdata = 32'd52747;
			12790: outdata = 32'd52746;
			12791: outdata = 32'd52745;
			12792: outdata = 32'd52744;
			12793: outdata = 32'd52743;
			12794: outdata = 32'd52742;
			12795: outdata = 32'd52741;
			12796: outdata = 32'd52740;
			12797: outdata = 32'd52739;
			12798: outdata = 32'd52738;
			12799: outdata = 32'd52737;
			12800: outdata = 32'd52736;
			12801: outdata = 32'd52735;
			12802: outdata = 32'd52734;
			12803: outdata = 32'd52733;
			12804: outdata = 32'd52732;
			12805: outdata = 32'd52731;
			12806: outdata = 32'd52730;
			12807: outdata = 32'd52729;
			12808: outdata = 32'd52728;
			12809: outdata = 32'd52727;
			12810: outdata = 32'd52726;
			12811: outdata = 32'd52725;
			12812: outdata = 32'd52724;
			12813: outdata = 32'd52723;
			12814: outdata = 32'd52722;
			12815: outdata = 32'd52721;
			12816: outdata = 32'd52720;
			12817: outdata = 32'd52719;
			12818: outdata = 32'd52718;
			12819: outdata = 32'd52717;
			12820: outdata = 32'd52716;
			12821: outdata = 32'd52715;
			12822: outdata = 32'd52714;
			12823: outdata = 32'd52713;
			12824: outdata = 32'd52712;
			12825: outdata = 32'd52711;
			12826: outdata = 32'd52710;
			12827: outdata = 32'd52709;
			12828: outdata = 32'd52708;
			12829: outdata = 32'd52707;
			12830: outdata = 32'd52706;
			12831: outdata = 32'd52705;
			12832: outdata = 32'd52704;
			12833: outdata = 32'd52703;
			12834: outdata = 32'd52702;
			12835: outdata = 32'd52701;
			12836: outdata = 32'd52700;
			12837: outdata = 32'd52699;
			12838: outdata = 32'd52698;
			12839: outdata = 32'd52697;
			12840: outdata = 32'd52696;
			12841: outdata = 32'd52695;
			12842: outdata = 32'd52694;
			12843: outdata = 32'd52693;
			12844: outdata = 32'd52692;
			12845: outdata = 32'd52691;
			12846: outdata = 32'd52690;
			12847: outdata = 32'd52689;
			12848: outdata = 32'd52688;
			12849: outdata = 32'd52687;
			12850: outdata = 32'd52686;
			12851: outdata = 32'd52685;
			12852: outdata = 32'd52684;
			12853: outdata = 32'd52683;
			12854: outdata = 32'd52682;
			12855: outdata = 32'd52681;
			12856: outdata = 32'd52680;
			12857: outdata = 32'd52679;
			12858: outdata = 32'd52678;
			12859: outdata = 32'd52677;
			12860: outdata = 32'd52676;
			12861: outdata = 32'd52675;
			12862: outdata = 32'd52674;
			12863: outdata = 32'd52673;
			12864: outdata = 32'd52672;
			12865: outdata = 32'd52671;
			12866: outdata = 32'd52670;
			12867: outdata = 32'd52669;
			12868: outdata = 32'd52668;
			12869: outdata = 32'd52667;
			12870: outdata = 32'd52666;
			12871: outdata = 32'd52665;
			12872: outdata = 32'd52664;
			12873: outdata = 32'd52663;
			12874: outdata = 32'd52662;
			12875: outdata = 32'd52661;
			12876: outdata = 32'd52660;
			12877: outdata = 32'd52659;
			12878: outdata = 32'd52658;
			12879: outdata = 32'd52657;
			12880: outdata = 32'd52656;
			12881: outdata = 32'd52655;
			12882: outdata = 32'd52654;
			12883: outdata = 32'd52653;
			12884: outdata = 32'd52652;
			12885: outdata = 32'd52651;
			12886: outdata = 32'd52650;
			12887: outdata = 32'd52649;
			12888: outdata = 32'd52648;
			12889: outdata = 32'd52647;
			12890: outdata = 32'd52646;
			12891: outdata = 32'd52645;
			12892: outdata = 32'd52644;
			12893: outdata = 32'd52643;
			12894: outdata = 32'd52642;
			12895: outdata = 32'd52641;
			12896: outdata = 32'd52640;
			12897: outdata = 32'd52639;
			12898: outdata = 32'd52638;
			12899: outdata = 32'd52637;
			12900: outdata = 32'd52636;
			12901: outdata = 32'd52635;
			12902: outdata = 32'd52634;
			12903: outdata = 32'd52633;
			12904: outdata = 32'd52632;
			12905: outdata = 32'd52631;
			12906: outdata = 32'd52630;
			12907: outdata = 32'd52629;
			12908: outdata = 32'd52628;
			12909: outdata = 32'd52627;
			12910: outdata = 32'd52626;
			12911: outdata = 32'd52625;
			12912: outdata = 32'd52624;
			12913: outdata = 32'd52623;
			12914: outdata = 32'd52622;
			12915: outdata = 32'd52621;
			12916: outdata = 32'd52620;
			12917: outdata = 32'd52619;
			12918: outdata = 32'd52618;
			12919: outdata = 32'd52617;
			12920: outdata = 32'd52616;
			12921: outdata = 32'd52615;
			12922: outdata = 32'd52614;
			12923: outdata = 32'd52613;
			12924: outdata = 32'd52612;
			12925: outdata = 32'd52611;
			12926: outdata = 32'd52610;
			12927: outdata = 32'd52609;
			12928: outdata = 32'd52608;
			12929: outdata = 32'd52607;
			12930: outdata = 32'd52606;
			12931: outdata = 32'd52605;
			12932: outdata = 32'd52604;
			12933: outdata = 32'd52603;
			12934: outdata = 32'd52602;
			12935: outdata = 32'd52601;
			12936: outdata = 32'd52600;
			12937: outdata = 32'd52599;
			12938: outdata = 32'd52598;
			12939: outdata = 32'd52597;
			12940: outdata = 32'd52596;
			12941: outdata = 32'd52595;
			12942: outdata = 32'd52594;
			12943: outdata = 32'd52593;
			12944: outdata = 32'd52592;
			12945: outdata = 32'd52591;
			12946: outdata = 32'd52590;
			12947: outdata = 32'd52589;
			12948: outdata = 32'd52588;
			12949: outdata = 32'd52587;
			12950: outdata = 32'd52586;
			12951: outdata = 32'd52585;
			12952: outdata = 32'd52584;
			12953: outdata = 32'd52583;
			12954: outdata = 32'd52582;
			12955: outdata = 32'd52581;
			12956: outdata = 32'd52580;
			12957: outdata = 32'd52579;
			12958: outdata = 32'd52578;
			12959: outdata = 32'd52577;
			12960: outdata = 32'd52576;
			12961: outdata = 32'd52575;
			12962: outdata = 32'd52574;
			12963: outdata = 32'd52573;
			12964: outdata = 32'd52572;
			12965: outdata = 32'd52571;
			12966: outdata = 32'd52570;
			12967: outdata = 32'd52569;
			12968: outdata = 32'd52568;
			12969: outdata = 32'd52567;
			12970: outdata = 32'd52566;
			12971: outdata = 32'd52565;
			12972: outdata = 32'd52564;
			12973: outdata = 32'd52563;
			12974: outdata = 32'd52562;
			12975: outdata = 32'd52561;
			12976: outdata = 32'd52560;
			12977: outdata = 32'd52559;
			12978: outdata = 32'd52558;
			12979: outdata = 32'd52557;
			12980: outdata = 32'd52556;
			12981: outdata = 32'd52555;
			12982: outdata = 32'd52554;
			12983: outdata = 32'd52553;
			12984: outdata = 32'd52552;
			12985: outdata = 32'd52551;
			12986: outdata = 32'd52550;
			12987: outdata = 32'd52549;
			12988: outdata = 32'd52548;
			12989: outdata = 32'd52547;
			12990: outdata = 32'd52546;
			12991: outdata = 32'd52545;
			12992: outdata = 32'd52544;
			12993: outdata = 32'd52543;
			12994: outdata = 32'd52542;
			12995: outdata = 32'd52541;
			12996: outdata = 32'd52540;
			12997: outdata = 32'd52539;
			12998: outdata = 32'd52538;
			12999: outdata = 32'd52537;
			13000: outdata = 32'd52536;
			13001: outdata = 32'd52535;
			13002: outdata = 32'd52534;
			13003: outdata = 32'd52533;
			13004: outdata = 32'd52532;
			13005: outdata = 32'd52531;
			13006: outdata = 32'd52530;
			13007: outdata = 32'd52529;
			13008: outdata = 32'd52528;
			13009: outdata = 32'd52527;
			13010: outdata = 32'd52526;
			13011: outdata = 32'd52525;
			13012: outdata = 32'd52524;
			13013: outdata = 32'd52523;
			13014: outdata = 32'd52522;
			13015: outdata = 32'd52521;
			13016: outdata = 32'd52520;
			13017: outdata = 32'd52519;
			13018: outdata = 32'd52518;
			13019: outdata = 32'd52517;
			13020: outdata = 32'd52516;
			13021: outdata = 32'd52515;
			13022: outdata = 32'd52514;
			13023: outdata = 32'd52513;
			13024: outdata = 32'd52512;
			13025: outdata = 32'd52511;
			13026: outdata = 32'd52510;
			13027: outdata = 32'd52509;
			13028: outdata = 32'd52508;
			13029: outdata = 32'd52507;
			13030: outdata = 32'd52506;
			13031: outdata = 32'd52505;
			13032: outdata = 32'd52504;
			13033: outdata = 32'd52503;
			13034: outdata = 32'd52502;
			13035: outdata = 32'd52501;
			13036: outdata = 32'd52500;
			13037: outdata = 32'd52499;
			13038: outdata = 32'd52498;
			13039: outdata = 32'd52497;
			13040: outdata = 32'd52496;
			13041: outdata = 32'd52495;
			13042: outdata = 32'd52494;
			13043: outdata = 32'd52493;
			13044: outdata = 32'd52492;
			13045: outdata = 32'd52491;
			13046: outdata = 32'd52490;
			13047: outdata = 32'd52489;
			13048: outdata = 32'd52488;
			13049: outdata = 32'd52487;
			13050: outdata = 32'd52486;
			13051: outdata = 32'd52485;
			13052: outdata = 32'd52484;
			13053: outdata = 32'd52483;
			13054: outdata = 32'd52482;
			13055: outdata = 32'd52481;
			13056: outdata = 32'd52480;
			13057: outdata = 32'd52479;
			13058: outdata = 32'd52478;
			13059: outdata = 32'd52477;
			13060: outdata = 32'd52476;
			13061: outdata = 32'd52475;
			13062: outdata = 32'd52474;
			13063: outdata = 32'd52473;
			13064: outdata = 32'd52472;
			13065: outdata = 32'd52471;
			13066: outdata = 32'd52470;
			13067: outdata = 32'd52469;
			13068: outdata = 32'd52468;
			13069: outdata = 32'd52467;
			13070: outdata = 32'd52466;
			13071: outdata = 32'd52465;
			13072: outdata = 32'd52464;
			13073: outdata = 32'd52463;
			13074: outdata = 32'd52462;
			13075: outdata = 32'd52461;
			13076: outdata = 32'd52460;
			13077: outdata = 32'd52459;
			13078: outdata = 32'd52458;
			13079: outdata = 32'd52457;
			13080: outdata = 32'd52456;
			13081: outdata = 32'd52455;
			13082: outdata = 32'd52454;
			13083: outdata = 32'd52453;
			13084: outdata = 32'd52452;
			13085: outdata = 32'd52451;
			13086: outdata = 32'd52450;
			13087: outdata = 32'd52449;
			13088: outdata = 32'd52448;
			13089: outdata = 32'd52447;
			13090: outdata = 32'd52446;
			13091: outdata = 32'd52445;
			13092: outdata = 32'd52444;
			13093: outdata = 32'd52443;
			13094: outdata = 32'd52442;
			13095: outdata = 32'd52441;
			13096: outdata = 32'd52440;
			13097: outdata = 32'd52439;
			13098: outdata = 32'd52438;
			13099: outdata = 32'd52437;
			13100: outdata = 32'd52436;
			13101: outdata = 32'd52435;
			13102: outdata = 32'd52434;
			13103: outdata = 32'd52433;
			13104: outdata = 32'd52432;
			13105: outdata = 32'd52431;
			13106: outdata = 32'd52430;
			13107: outdata = 32'd52429;
			13108: outdata = 32'd52428;
			13109: outdata = 32'd52427;
			13110: outdata = 32'd52426;
			13111: outdata = 32'd52425;
			13112: outdata = 32'd52424;
			13113: outdata = 32'd52423;
			13114: outdata = 32'd52422;
			13115: outdata = 32'd52421;
			13116: outdata = 32'd52420;
			13117: outdata = 32'd52419;
			13118: outdata = 32'd52418;
			13119: outdata = 32'd52417;
			13120: outdata = 32'd52416;
			13121: outdata = 32'd52415;
			13122: outdata = 32'd52414;
			13123: outdata = 32'd52413;
			13124: outdata = 32'd52412;
			13125: outdata = 32'd52411;
			13126: outdata = 32'd52410;
			13127: outdata = 32'd52409;
			13128: outdata = 32'd52408;
			13129: outdata = 32'd52407;
			13130: outdata = 32'd52406;
			13131: outdata = 32'd52405;
			13132: outdata = 32'd52404;
			13133: outdata = 32'd52403;
			13134: outdata = 32'd52402;
			13135: outdata = 32'd52401;
			13136: outdata = 32'd52400;
			13137: outdata = 32'd52399;
			13138: outdata = 32'd52398;
			13139: outdata = 32'd52397;
			13140: outdata = 32'd52396;
			13141: outdata = 32'd52395;
			13142: outdata = 32'd52394;
			13143: outdata = 32'd52393;
			13144: outdata = 32'd52392;
			13145: outdata = 32'd52391;
			13146: outdata = 32'd52390;
			13147: outdata = 32'd52389;
			13148: outdata = 32'd52388;
			13149: outdata = 32'd52387;
			13150: outdata = 32'd52386;
			13151: outdata = 32'd52385;
			13152: outdata = 32'd52384;
			13153: outdata = 32'd52383;
			13154: outdata = 32'd52382;
			13155: outdata = 32'd52381;
			13156: outdata = 32'd52380;
			13157: outdata = 32'd52379;
			13158: outdata = 32'd52378;
			13159: outdata = 32'd52377;
			13160: outdata = 32'd52376;
			13161: outdata = 32'd52375;
			13162: outdata = 32'd52374;
			13163: outdata = 32'd52373;
			13164: outdata = 32'd52372;
			13165: outdata = 32'd52371;
			13166: outdata = 32'd52370;
			13167: outdata = 32'd52369;
			13168: outdata = 32'd52368;
			13169: outdata = 32'd52367;
			13170: outdata = 32'd52366;
			13171: outdata = 32'd52365;
			13172: outdata = 32'd52364;
			13173: outdata = 32'd52363;
			13174: outdata = 32'd52362;
			13175: outdata = 32'd52361;
			13176: outdata = 32'd52360;
			13177: outdata = 32'd52359;
			13178: outdata = 32'd52358;
			13179: outdata = 32'd52357;
			13180: outdata = 32'd52356;
			13181: outdata = 32'd52355;
			13182: outdata = 32'd52354;
			13183: outdata = 32'd52353;
			13184: outdata = 32'd52352;
			13185: outdata = 32'd52351;
			13186: outdata = 32'd52350;
			13187: outdata = 32'd52349;
			13188: outdata = 32'd52348;
			13189: outdata = 32'd52347;
			13190: outdata = 32'd52346;
			13191: outdata = 32'd52345;
			13192: outdata = 32'd52344;
			13193: outdata = 32'd52343;
			13194: outdata = 32'd52342;
			13195: outdata = 32'd52341;
			13196: outdata = 32'd52340;
			13197: outdata = 32'd52339;
			13198: outdata = 32'd52338;
			13199: outdata = 32'd52337;
			13200: outdata = 32'd52336;
			13201: outdata = 32'd52335;
			13202: outdata = 32'd52334;
			13203: outdata = 32'd52333;
			13204: outdata = 32'd52332;
			13205: outdata = 32'd52331;
			13206: outdata = 32'd52330;
			13207: outdata = 32'd52329;
			13208: outdata = 32'd52328;
			13209: outdata = 32'd52327;
			13210: outdata = 32'd52326;
			13211: outdata = 32'd52325;
			13212: outdata = 32'd52324;
			13213: outdata = 32'd52323;
			13214: outdata = 32'd52322;
			13215: outdata = 32'd52321;
			13216: outdata = 32'd52320;
			13217: outdata = 32'd52319;
			13218: outdata = 32'd52318;
			13219: outdata = 32'd52317;
			13220: outdata = 32'd52316;
			13221: outdata = 32'd52315;
			13222: outdata = 32'd52314;
			13223: outdata = 32'd52313;
			13224: outdata = 32'd52312;
			13225: outdata = 32'd52311;
			13226: outdata = 32'd52310;
			13227: outdata = 32'd52309;
			13228: outdata = 32'd52308;
			13229: outdata = 32'd52307;
			13230: outdata = 32'd52306;
			13231: outdata = 32'd52305;
			13232: outdata = 32'd52304;
			13233: outdata = 32'd52303;
			13234: outdata = 32'd52302;
			13235: outdata = 32'd52301;
			13236: outdata = 32'd52300;
			13237: outdata = 32'd52299;
			13238: outdata = 32'd52298;
			13239: outdata = 32'd52297;
			13240: outdata = 32'd52296;
			13241: outdata = 32'd52295;
			13242: outdata = 32'd52294;
			13243: outdata = 32'd52293;
			13244: outdata = 32'd52292;
			13245: outdata = 32'd52291;
			13246: outdata = 32'd52290;
			13247: outdata = 32'd52289;
			13248: outdata = 32'd52288;
			13249: outdata = 32'd52287;
			13250: outdata = 32'd52286;
			13251: outdata = 32'd52285;
			13252: outdata = 32'd52284;
			13253: outdata = 32'd52283;
			13254: outdata = 32'd52282;
			13255: outdata = 32'd52281;
			13256: outdata = 32'd52280;
			13257: outdata = 32'd52279;
			13258: outdata = 32'd52278;
			13259: outdata = 32'd52277;
			13260: outdata = 32'd52276;
			13261: outdata = 32'd52275;
			13262: outdata = 32'd52274;
			13263: outdata = 32'd52273;
			13264: outdata = 32'd52272;
			13265: outdata = 32'd52271;
			13266: outdata = 32'd52270;
			13267: outdata = 32'd52269;
			13268: outdata = 32'd52268;
			13269: outdata = 32'd52267;
			13270: outdata = 32'd52266;
			13271: outdata = 32'd52265;
			13272: outdata = 32'd52264;
			13273: outdata = 32'd52263;
			13274: outdata = 32'd52262;
			13275: outdata = 32'd52261;
			13276: outdata = 32'd52260;
			13277: outdata = 32'd52259;
			13278: outdata = 32'd52258;
			13279: outdata = 32'd52257;
			13280: outdata = 32'd52256;
			13281: outdata = 32'd52255;
			13282: outdata = 32'd52254;
			13283: outdata = 32'd52253;
			13284: outdata = 32'd52252;
			13285: outdata = 32'd52251;
			13286: outdata = 32'd52250;
			13287: outdata = 32'd52249;
			13288: outdata = 32'd52248;
			13289: outdata = 32'd52247;
			13290: outdata = 32'd52246;
			13291: outdata = 32'd52245;
			13292: outdata = 32'd52244;
			13293: outdata = 32'd52243;
			13294: outdata = 32'd52242;
			13295: outdata = 32'd52241;
			13296: outdata = 32'd52240;
			13297: outdata = 32'd52239;
			13298: outdata = 32'd52238;
			13299: outdata = 32'd52237;
			13300: outdata = 32'd52236;
			13301: outdata = 32'd52235;
			13302: outdata = 32'd52234;
			13303: outdata = 32'd52233;
			13304: outdata = 32'd52232;
			13305: outdata = 32'd52231;
			13306: outdata = 32'd52230;
			13307: outdata = 32'd52229;
			13308: outdata = 32'd52228;
			13309: outdata = 32'd52227;
			13310: outdata = 32'd52226;
			13311: outdata = 32'd52225;
			13312: outdata = 32'd52224;
			13313: outdata = 32'd52223;
			13314: outdata = 32'd52222;
			13315: outdata = 32'd52221;
			13316: outdata = 32'd52220;
			13317: outdata = 32'd52219;
			13318: outdata = 32'd52218;
			13319: outdata = 32'd52217;
			13320: outdata = 32'd52216;
			13321: outdata = 32'd52215;
			13322: outdata = 32'd52214;
			13323: outdata = 32'd52213;
			13324: outdata = 32'd52212;
			13325: outdata = 32'd52211;
			13326: outdata = 32'd52210;
			13327: outdata = 32'd52209;
			13328: outdata = 32'd52208;
			13329: outdata = 32'd52207;
			13330: outdata = 32'd52206;
			13331: outdata = 32'd52205;
			13332: outdata = 32'd52204;
			13333: outdata = 32'd52203;
			13334: outdata = 32'd52202;
			13335: outdata = 32'd52201;
			13336: outdata = 32'd52200;
			13337: outdata = 32'd52199;
			13338: outdata = 32'd52198;
			13339: outdata = 32'd52197;
			13340: outdata = 32'd52196;
			13341: outdata = 32'd52195;
			13342: outdata = 32'd52194;
			13343: outdata = 32'd52193;
			13344: outdata = 32'd52192;
			13345: outdata = 32'd52191;
			13346: outdata = 32'd52190;
			13347: outdata = 32'd52189;
			13348: outdata = 32'd52188;
			13349: outdata = 32'd52187;
			13350: outdata = 32'd52186;
			13351: outdata = 32'd52185;
			13352: outdata = 32'd52184;
			13353: outdata = 32'd52183;
			13354: outdata = 32'd52182;
			13355: outdata = 32'd52181;
			13356: outdata = 32'd52180;
			13357: outdata = 32'd52179;
			13358: outdata = 32'd52178;
			13359: outdata = 32'd52177;
			13360: outdata = 32'd52176;
			13361: outdata = 32'd52175;
			13362: outdata = 32'd52174;
			13363: outdata = 32'd52173;
			13364: outdata = 32'd52172;
			13365: outdata = 32'd52171;
			13366: outdata = 32'd52170;
			13367: outdata = 32'd52169;
			13368: outdata = 32'd52168;
			13369: outdata = 32'd52167;
			13370: outdata = 32'd52166;
			13371: outdata = 32'd52165;
			13372: outdata = 32'd52164;
			13373: outdata = 32'd52163;
			13374: outdata = 32'd52162;
			13375: outdata = 32'd52161;
			13376: outdata = 32'd52160;
			13377: outdata = 32'd52159;
			13378: outdata = 32'd52158;
			13379: outdata = 32'd52157;
			13380: outdata = 32'd52156;
			13381: outdata = 32'd52155;
			13382: outdata = 32'd52154;
			13383: outdata = 32'd52153;
			13384: outdata = 32'd52152;
			13385: outdata = 32'd52151;
			13386: outdata = 32'd52150;
			13387: outdata = 32'd52149;
			13388: outdata = 32'd52148;
			13389: outdata = 32'd52147;
			13390: outdata = 32'd52146;
			13391: outdata = 32'd52145;
			13392: outdata = 32'd52144;
			13393: outdata = 32'd52143;
			13394: outdata = 32'd52142;
			13395: outdata = 32'd52141;
			13396: outdata = 32'd52140;
			13397: outdata = 32'd52139;
			13398: outdata = 32'd52138;
			13399: outdata = 32'd52137;
			13400: outdata = 32'd52136;
			13401: outdata = 32'd52135;
			13402: outdata = 32'd52134;
			13403: outdata = 32'd52133;
			13404: outdata = 32'd52132;
			13405: outdata = 32'd52131;
			13406: outdata = 32'd52130;
			13407: outdata = 32'd52129;
			13408: outdata = 32'd52128;
			13409: outdata = 32'd52127;
			13410: outdata = 32'd52126;
			13411: outdata = 32'd52125;
			13412: outdata = 32'd52124;
			13413: outdata = 32'd52123;
			13414: outdata = 32'd52122;
			13415: outdata = 32'd52121;
			13416: outdata = 32'd52120;
			13417: outdata = 32'd52119;
			13418: outdata = 32'd52118;
			13419: outdata = 32'd52117;
			13420: outdata = 32'd52116;
			13421: outdata = 32'd52115;
			13422: outdata = 32'd52114;
			13423: outdata = 32'd52113;
			13424: outdata = 32'd52112;
			13425: outdata = 32'd52111;
			13426: outdata = 32'd52110;
			13427: outdata = 32'd52109;
			13428: outdata = 32'd52108;
			13429: outdata = 32'd52107;
			13430: outdata = 32'd52106;
			13431: outdata = 32'd52105;
			13432: outdata = 32'd52104;
			13433: outdata = 32'd52103;
			13434: outdata = 32'd52102;
			13435: outdata = 32'd52101;
			13436: outdata = 32'd52100;
			13437: outdata = 32'd52099;
			13438: outdata = 32'd52098;
			13439: outdata = 32'd52097;
			13440: outdata = 32'd52096;
			13441: outdata = 32'd52095;
			13442: outdata = 32'd52094;
			13443: outdata = 32'd52093;
			13444: outdata = 32'd52092;
			13445: outdata = 32'd52091;
			13446: outdata = 32'd52090;
			13447: outdata = 32'd52089;
			13448: outdata = 32'd52088;
			13449: outdata = 32'd52087;
			13450: outdata = 32'd52086;
			13451: outdata = 32'd52085;
			13452: outdata = 32'd52084;
			13453: outdata = 32'd52083;
			13454: outdata = 32'd52082;
			13455: outdata = 32'd52081;
			13456: outdata = 32'd52080;
			13457: outdata = 32'd52079;
			13458: outdata = 32'd52078;
			13459: outdata = 32'd52077;
			13460: outdata = 32'd52076;
			13461: outdata = 32'd52075;
			13462: outdata = 32'd52074;
			13463: outdata = 32'd52073;
			13464: outdata = 32'd52072;
			13465: outdata = 32'd52071;
			13466: outdata = 32'd52070;
			13467: outdata = 32'd52069;
			13468: outdata = 32'd52068;
			13469: outdata = 32'd52067;
			13470: outdata = 32'd52066;
			13471: outdata = 32'd52065;
			13472: outdata = 32'd52064;
			13473: outdata = 32'd52063;
			13474: outdata = 32'd52062;
			13475: outdata = 32'd52061;
			13476: outdata = 32'd52060;
			13477: outdata = 32'd52059;
			13478: outdata = 32'd52058;
			13479: outdata = 32'd52057;
			13480: outdata = 32'd52056;
			13481: outdata = 32'd52055;
			13482: outdata = 32'd52054;
			13483: outdata = 32'd52053;
			13484: outdata = 32'd52052;
			13485: outdata = 32'd52051;
			13486: outdata = 32'd52050;
			13487: outdata = 32'd52049;
			13488: outdata = 32'd52048;
			13489: outdata = 32'd52047;
			13490: outdata = 32'd52046;
			13491: outdata = 32'd52045;
			13492: outdata = 32'd52044;
			13493: outdata = 32'd52043;
			13494: outdata = 32'd52042;
			13495: outdata = 32'd52041;
			13496: outdata = 32'd52040;
			13497: outdata = 32'd52039;
			13498: outdata = 32'd52038;
			13499: outdata = 32'd52037;
			13500: outdata = 32'd52036;
			13501: outdata = 32'd52035;
			13502: outdata = 32'd52034;
			13503: outdata = 32'd52033;
			13504: outdata = 32'd52032;
			13505: outdata = 32'd52031;
			13506: outdata = 32'd52030;
			13507: outdata = 32'd52029;
			13508: outdata = 32'd52028;
			13509: outdata = 32'd52027;
			13510: outdata = 32'd52026;
			13511: outdata = 32'd52025;
			13512: outdata = 32'd52024;
			13513: outdata = 32'd52023;
			13514: outdata = 32'd52022;
			13515: outdata = 32'd52021;
			13516: outdata = 32'd52020;
			13517: outdata = 32'd52019;
			13518: outdata = 32'd52018;
			13519: outdata = 32'd52017;
			13520: outdata = 32'd52016;
			13521: outdata = 32'd52015;
			13522: outdata = 32'd52014;
			13523: outdata = 32'd52013;
			13524: outdata = 32'd52012;
			13525: outdata = 32'd52011;
			13526: outdata = 32'd52010;
			13527: outdata = 32'd52009;
			13528: outdata = 32'd52008;
			13529: outdata = 32'd52007;
			13530: outdata = 32'd52006;
			13531: outdata = 32'd52005;
			13532: outdata = 32'd52004;
			13533: outdata = 32'd52003;
			13534: outdata = 32'd52002;
			13535: outdata = 32'd52001;
			13536: outdata = 32'd52000;
			13537: outdata = 32'd51999;
			13538: outdata = 32'd51998;
			13539: outdata = 32'd51997;
			13540: outdata = 32'd51996;
			13541: outdata = 32'd51995;
			13542: outdata = 32'd51994;
			13543: outdata = 32'd51993;
			13544: outdata = 32'd51992;
			13545: outdata = 32'd51991;
			13546: outdata = 32'd51990;
			13547: outdata = 32'd51989;
			13548: outdata = 32'd51988;
			13549: outdata = 32'd51987;
			13550: outdata = 32'd51986;
			13551: outdata = 32'd51985;
			13552: outdata = 32'd51984;
			13553: outdata = 32'd51983;
			13554: outdata = 32'd51982;
			13555: outdata = 32'd51981;
			13556: outdata = 32'd51980;
			13557: outdata = 32'd51979;
			13558: outdata = 32'd51978;
			13559: outdata = 32'd51977;
			13560: outdata = 32'd51976;
			13561: outdata = 32'd51975;
			13562: outdata = 32'd51974;
			13563: outdata = 32'd51973;
			13564: outdata = 32'd51972;
			13565: outdata = 32'd51971;
			13566: outdata = 32'd51970;
			13567: outdata = 32'd51969;
			13568: outdata = 32'd51968;
			13569: outdata = 32'd51967;
			13570: outdata = 32'd51966;
			13571: outdata = 32'd51965;
			13572: outdata = 32'd51964;
			13573: outdata = 32'd51963;
			13574: outdata = 32'd51962;
			13575: outdata = 32'd51961;
			13576: outdata = 32'd51960;
			13577: outdata = 32'd51959;
			13578: outdata = 32'd51958;
			13579: outdata = 32'd51957;
			13580: outdata = 32'd51956;
			13581: outdata = 32'd51955;
			13582: outdata = 32'd51954;
			13583: outdata = 32'd51953;
			13584: outdata = 32'd51952;
			13585: outdata = 32'd51951;
			13586: outdata = 32'd51950;
			13587: outdata = 32'd51949;
			13588: outdata = 32'd51948;
			13589: outdata = 32'd51947;
			13590: outdata = 32'd51946;
			13591: outdata = 32'd51945;
			13592: outdata = 32'd51944;
			13593: outdata = 32'd51943;
			13594: outdata = 32'd51942;
			13595: outdata = 32'd51941;
			13596: outdata = 32'd51940;
			13597: outdata = 32'd51939;
			13598: outdata = 32'd51938;
			13599: outdata = 32'd51937;
			13600: outdata = 32'd51936;
			13601: outdata = 32'd51935;
			13602: outdata = 32'd51934;
			13603: outdata = 32'd51933;
			13604: outdata = 32'd51932;
			13605: outdata = 32'd51931;
			13606: outdata = 32'd51930;
			13607: outdata = 32'd51929;
			13608: outdata = 32'd51928;
			13609: outdata = 32'd51927;
			13610: outdata = 32'd51926;
			13611: outdata = 32'd51925;
			13612: outdata = 32'd51924;
			13613: outdata = 32'd51923;
			13614: outdata = 32'd51922;
			13615: outdata = 32'd51921;
			13616: outdata = 32'd51920;
			13617: outdata = 32'd51919;
			13618: outdata = 32'd51918;
			13619: outdata = 32'd51917;
			13620: outdata = 32'd51916;
			13621: outdata = 32'd51915;
			13622: outdata = 32'd51914;
			13623: outdata = 32'd51913;
			13624: outdata = 32'd51912;
			13625: outdata = 32'd51911;
			13626: outdata = 32'd51910;
			13627: outdata = 32'd51909;
			13628: outdata = 32'd51908;
			13629: outdata = 32'd51907;
			13630: outdata = 32'd51906;
			13631: outdata = 32'd51905;
			13632: outdata = 32'd51904;
			13633: outdata = 32'd51903;
			13634: outdata = 32'd51902;
			13635: outdata = 32'd51901;
			13636: outdata = 32'd51900;
			13637: outdata = 32'd51899;
			13638: outdata = 32'd51898;
			13639: outdata = 32'd51897;
			13640: outdata = 32'd51896;
			13641: outdata = 32'd51895;
			13642: outdata = 32'd51894;
			13643: outdata = 32'd51893;
			13644: outdata = 32'd51892;
			13645: outdata = 32'd51891;
			13646: outdata = 32'd51890;
			13647: outdata = 32'd51889;
			13648: outdata = 32'd51888;
			13649: outdata = 32'd51887;
			13650: outdata = 32'd51886;
			13651: outdata = 32'd51885;
			13652: outdata = 32'd51884;
			13653: outdata = 32'd51883;
			13654: outdata = 32'd51882;
			13655: outdata = 32'd51881;
			13656: outdata = 32'd51880;
			13657: outdata = 32'd51879;
			13658: outdata = 32'd51878;
			13659: outdata = 32'd51877;
			13660: outdata = 32'd51876;
			13661: outdata = 32'd51875;
			13662: outdata = 32'd51874;
			13663: outdata = 32'd51873;
			13664: outdata = 32'd51872;
			13665: outdata = 32'd51871;
			13666: outdata = 32'd51870;
			13667: outdata = 32'd51869;
			13668: outdata = 32'd51868;
			13669: outdata = 32'd51867;
			13670: outdata = 32'd51866;
			13671: outdata = 32'd51865;
			13672: outdata = 32'd51864;
			13673: outdata = 32'd51863;
			13674: outdata = 32'd51862;
			13675: outdata = 32'd51861;
			13676: outdata = 32'd51860;
			13677: outdata = 32'd51859;
			13678: outdata = 32'd51858;
			13679: outdata = 32'd51857;
			13680: outdata = 32'd51856;
			13681: outdata = 32'd51855;
			13682: outdata = 32'd51854;
			13683: outdata = 32'd51853;
			13684: outdata = 32'd51852;
			13685: outdata = 32'd51851;
			13686: outdata = 32'd51850;
			13687: outdata = 32'd51849;
			13688: outdata = 32'd51848;
			13689: outdata = 32'd51847;
			13690: outdata = 32'd51846;
			13691: outdata = 32'd51845;
			13692: outdata = 32'd51844;
			13693: outdata = 32'd51843;
			13694: outdata = 32'd51842;
			13695: outdata = 32'd51841;
			13696: outdata = 32'd51840;
			13697: outdata = 32'd51839;
			13698: outdata = 32'd51838;
			13699: outdata = 32'd51837;
			13700: outdata = 32'd51836;
			13701: outdata = 32'd51835;
			13702: outdata = 32'd51834;
			13703: outdata = 32'd51833;
			13704: outdata = 32'd51832;
			13705: outdata = 32'd51831;
			13706: outdata = 32'd51830;
			13707: outdata = 32'd51829;
			13708: outdata = 32'd51828;
			13709: outdata = 32'd51827;
			13710: outdata = 32'd51826;
			13711: outdata = 32'd51825;
			13712: outdata = 32'd51824;
			13713: outdata = 32'd51823;
			13714: outdata = 32'd51822;
			13715: outdata = 32'd51821;
			13716: outdata = 32'd51820;
			13717: outdata = 32'd51819;
			13718: outdata = 32'd51818;
			13719: outdata = 32'd51817;
			13720: outdata = 32'd51816;
			13721: outdata = 32'd51815;
			13722: outdata = 32'd51814;
			13723: outdata = 32'd51813;
			13724: outdata = 32'd51812;
			13725: outdata = 32'd51811;
			13726: outdata = 32'd51810;
			13727: outdata = 32'd51809;
			13728: outdata = 32'd51808;
			13729: outdata = 32'd51807;
			13730: outdata = 32'd51806;
			13731: outdata = 32'd51805;
			13732: outdata = 32'd51804;
			13733: outdata = 32'd51803;
			13734: outdata = 32'd51802;
			13735: outdata = 32'd51801;
			13736: outdata = 32'd51800;
			13737: outdata = 32'd51799;
			13738: outdata = 32'd51798;
			13739: outdata = 32'd51797;
			13740: outdata = 32'd51796;
			13741: outdata = 32'd51795;
			13742: outdata = 32'd51794;
			13743: outdata = 32'd51793;
			13744: outdata = 32'd51792;
			13745: outdata = 32'd51791;
			13746: outdata = 32'd51790;
			13747: outdata = 32'd51789;
			13748: outdata = 32'd51788;
			13749: outdata = 32'd51787;
			13750: outdata = 32'd51786;
			13751: outdata = 32'd51785;
			13752: outdata = 32'd51784;
			13753: outdata = 32'd51783;
			13754: outdata = 32'd51782;
			13755: outdata = 32'd51781;
			13756: outdata = 32'd51780;
			13757: outdata = 32'd51779;
			13758: outdata = 32'd51778;
			13759: outdata = 32'd51777;
			13760: outdata = 32'd51776;
			13761: outdata = 32'd51775;
			13762: outdata = 32'd51774;
			13763: outdata = 32'd51773;
			13764: outdata = 32'd51772;
			13765: outdata = 32'd51771;
			13766: outdata = 32'd51770;
			13767: outdata = 32'd51769;
			13768: outdata = 32'd51768;
			13769: outdata = 32'd51767;
			13770: outdata = 32'd51766;
			13771: outdata = 32'd51765;
			13772: outdata = 32'd51764;
			13773: outdata = 32'd51763;
			13774: outdata = 32'd51762;
			13775: outdata = 32'd51761;
			13776: outdata = 32'd51760;
			13777: outdata = 32'd51759;
			13778: outdata = 32'd51758;
			13779: outdata = 32'd51757;
			13780: outdata = 32'd51756;
			13781: outdata = 32'd51755;
			13782: outdata = 32'd51754;
			13783: outdata = 32'd51753;
			13784: outdata = 32'd51752;
			13785: outdata = 32'd51751;
			13786: outdata = 32'd51750;
			13787: outdata = 32'd51749;
			13788: outdata = 32'd51748;
			13789: outdata = 32'd51747;
			13790: outdata = 32'd51746;
			13791: outdata = 32'd51745;
			13792: outdata = 32'd51744;
			13793: outdata = 32'd51743;
			13794: outdata = 32'd51742;
			13795: outdata = 32'd51741;
			13796: outdata = 32'd51740;
			13797: outdata = 32'd51739;
			13798: outdata = 32'd51738;
			13799: outdata = 32'd51737;
			13800: outdata = 32'd51736;
			13801: outdata = 32'd51735;
			13802: outdata = 32'd51734;
			13803: outdata = 32'd51733;
			13804: outdata = 32'd51732;
			13805: outdata = 32'd51731;
			13806: outdata = 32'd51730;
			13807: outdata = 32'd51729;
			13808: outdata = 32'd51728;
			13809: outdata = 32'd51727;
			13810: outdata = 32'd51726;
			13811: outdata = 32'd51725;
			13812: outdata = 32'd51724;
			13813: outdata = 32'd51723;
			13814: outdata = 32'd51722;
			13815: outdata = 32'd51721;
			13816: outdata = 32'd51720;
			13817: outdata = 32'd51719;
			13818: outdata = 32'd51718;
			13819: outdata = 32'd51717;
			13820: outdata = 32'd51716;
			13821: outdata = 32'd51715;
			13822: outdata = 32'd51714;
			13823: outdata = 32'd51713;
			13824: outdata = 32'd51712;
			13825: outdata = 32'd51711;
			13826: outdata = 32'd51710;
			13827: outdata = 32'd51709;
			13828: outdata = 32'd51708;
			13829: outdata = 32'd51707;
			13830: outdata = 32'd51706;
			13831: outdata = 32'd51705;
			13832: outdata = 32'd51704;
			13833: outdata = 32'd51703;
			13834: outdata = 32'd51702;
			13835: outdata = 32'd51701;
			13836: outdata = 32'd51700;
			13837: outdata = 32'd51699;
			13838: outdata = 32'd51698;
			13839: outdata = 32'd51697;
			13840: outdata = 32'd51696;
			13841: outdata = 32'd51695;
			13842: outdata = 32'd51694;
			13843: outdata = 32'd51693;
			13844: outdata = 32'd51692;
			13845: outdata = 32'd51691;
			13846: outdata = 32'd51690;
			13847: outdata = 32'd51689;
			13848: outdata = 32'd51688;
			13849: outdata = 32'd51687;
			13850: outdata = 32'd51686;
			13851: outdata = 32'd51685;
			13852: outdata = 32'd51684;
			13853: outdata = 32'd51683;
			13854: outdata = 32'd51682;
			13855: outdata = 32'd51681;
			13856: outdata = 32'd51680;
			13857: outdata = 32'd51679;
			13858: outdata = 32'd51678;
			13859: outdata = 32'd51677;
			13860: outdata = 32'd51676;
			13861: outdata = 32'd51675;
			13862: outdata = 32'd51674;
			13863: outdata = 32'd51673;
			13864: outdata = 32'd51672;
			13865: outdata = 32'd51671;
			13866: outdata = 32'd51670;
			13867: outdata = 32'd51669;
			13868: outdata = 32'd51668;
			13869: outdata = 32'd51667;
			13870: outdata = 32'd51666;
			13871: outdata = 32'd51665;
			13872: outdata = 32'd51664;
			13873: outdata = 32'd51663;
			13874: outdata = 32'd51662;
			13875: outdata = 32'd51661;
			13876: outdata = 32'd51660;
			13877: outdata = 32'd51659;
			13878: outdata = 32'd51658;
			13879: outdata = 32'd51657;
			13880: outdata = 32'd51656;
			13881: outdata = 32'd51655;
			13882: outdata = 32'd51654;
			13883: outdata = 32'd51653;
			13884: outdata = 32'd51652;
			13885: outdata = 32'd51651;
			13886: outdata = 32'd51650;
			13887: outdata = 32'd51649;
			13888: outdata = 32'd51648;
			13889: outdata = 32'd51647;
			13890: outdata = 32'd51646;
			13891: outdata = 32'd51645;
			13892: outdata = 32'd51644;
			13893: outdata = 32'd51643;
			13894: outdata = 32'd51642;
			13895: outdata = 32'd51641;
			13896: outdata = 32'd51640;
			13897: outdata = 32'd51639;
			13898: outdata = 32'd51638;
			13899: outdata = 32'd51637;
			13900: outdata = 32'd51636;
			13901: outdata = 32'd51635;
			13902: outdata = 32'd51634;
			13903: outdata = 32'd51633;
			13904: outdata = 32'd51632;
			13905: outdata = 32'd51631;
			13906: outdata = 32'd51630;
			13907: outdata = 32'd51629;
			13908: outdata = 32'd51628;
			13909: outdata = 32'd51627;
			13910: outdata = 32'd51626;
			13911: outdata = 32'd51625;
			13912: outdata = 32'd51624;
			13913: outdata = 32'd51623;
			13914: outdata = 32'd51622;
			13915: outdata = 32'd51621;
			13916: outdata = 32'd51620;
			13917: outdata = 32'd51619;
			13918: outdata = 32'd51618;
			13919: outdata = 32'd51617;
			13920: outdata = 32'd51616;
			13921: outdata = 32'd51615;
			13922: outdata = 32'd51614;
			13923: outdata = 32'd51613;
			13924: outdata = 32'd51612;
			13925: outdata = 32'd51611;
			13926: outdata = 32'd51610;
			13927: outdata = 32'd51609;
			13928: outdata = 32'd51608;
			13929: outdata = 32'd51607;
			13930: outdata = 32'd51606;
			13931: outdata = 32'd51605;
			13932: outdata = 32'd51604;
			13933: outdata = 32'd51603;
			13934: outdata = 32'd51602;
			13935: outdata = 32'd51601;
			13936: outdata = 32'd51600;
			13937: outdata = 32'd51599;
			13938: outdata = 32'd51598;
			13939: outdata = 32'd51597;
			13940: outdata = 32'd51596;
			13941: outdata = 32'd51595;
			13942: outdata = 32'd51594;
			13943: outdata = 32'd51593;
			13944: outdata = 32'd51592;
			13945: outdata = 32'd51591;
			13946: outdata = 32'd51590;
			13947: outdata = 32'd51589;
			13948: outdata = 32'd51588;
			13949: outdata = 32'd51587;
			13950: outdata = 32'd51586;
			13951: outdata = 32'd51585;
			13952: outdata = 32'd51584;
			13953: outdata = 32'd51583;
			13954: outdata = 32'd51582;
			13955: outdata = 32'd51581;
			13956: outdata = 32'd51580;
			13957: outdata = 32'd51579;
			13958: outdata = 32'd51578;
			13959: outdata = 32'd51577;
			13960: outdata = 32'd51576;
			13961: outdata = 32'd51575;
			13962: outdata = 32'd51574;
			13963: outdata = 32'd51573;
			13964: outdata = 32'd51572;
			13965: outdata = 32'd51571;
			13966: outdata = 32'd51570;
			13967: outdata = 32'd51569;
			13968: outdata = 32'd51568;
			13969: outdata = 32'd51567;
			13970: outdata = 32'd51566;
			13971: outdata = 32'd51565;
			13972: outdata = 32'd51564;
			13973: outdata = 32'd51563;
			13974: outdata = 32'd51562;
			13975: outdata = 32'd51561;
			13976: outdata = 32'd51560;
			13977: outdata = 32'd51559;
			13978: outdata = 32'd51558;
			13979: outdata = 32'd51557;
			13980: outdata = 32'd51556;
			13981: outdata = 32'd51555;
			13982: outdata = 32'd51554;
			13983: outdata = 32'd51553;
			13984: outdata = 32'd51552;
			13985: outdata = 32'd51551;
			13986: outdata = 32'd51550;
			13987: outdata = 32'd51549;
			13988: outdata = 32'd51548;
			13989: outdata = 32'd51547;
			13990: outdata = 32'd51546;
			13991: outdata = 32'd51545;
			13992: outdata = 32'd51544;
			13993: outdata = 32'd51543;
			13994: outdata = 32'd51542;
			13995: outdata = 32'd51541;
			13996: outdata = 32'd51540;
			13997: outdata = 32'd51539;
			13998: outdata = 32'd51538;
			13999: outdata = 32'd51537;
			14000: outdata = 32'd51536;
			14001: outdata = 32'd51535;
			14002: outdata = 32'd51534;
			14003: outdata = 32'd51533;
			14004: outdata = 32'd51532;
			14005: outdata = 32'd51531;
			14006: outdata = 32'd51530;
			14007: outdata = 32'd51529;
			14008: outdata = 32'd51528;
			14009: outdata = 32'd51527;
			14010: outdata = 32'd51526;
			14011: outdata = 32'd51525;
			14012: outdata = 32'd51524;
			14013: outdata = 32'd51523;
			14014: outdata = 32'd51522;
			14015: outdata = 32'd51521;
			14016: outdata = 32'd51520;
			14017: outdata = 32'd51519;
			14018: outdata = 32'd51518;
			14019: outdata = 32'd51517;
			14020: outdata = 32'd51516;
			14021: outdata = 32'd51515;
			14022: outdata = 32'd51514;
			14023: outdata = 32'd51513;
			14024: outdata = 32'd51512;
			14025: outdata = 32'd51511;
			14026: outdata = 32'd51510;
			14027: outdata = 32'd51509;
			14028: outdata = 32'd51508;
			14029: outdata = 32'd51507;
			14030: outdata = 32'd51506;
			14031: outdata = 32'd51505;
			14032: outdata = 32'd51504;
			14033: outdata = 32'd51503;
			14034: outdata = 32'd51502;
			14035: outdata = 32'd51501;
			14036: outdata = 32'd51500;
			14037: outdata = 32'd51499;
			14038: outdata = 32'd51498;
			14039: outdata = 32'd51497;
			14040: outdata = 32'd51496;
			14041: outdata = 32'd51495;
			14042: outdata = 32'd51494;
			14043: outdata = 32'd51493;
			14044: outdata = 32'd51492;
			14045: outdata = 32'd51491;
			14046: outdata = 32'd51490;
			14047: outdata = 32'd51489;
			14048: outdata = 32'd51488;
			14049: outdata = 32'd51487;
			14050: outdata = 32'd51486;
			14051: outdata = 32'd51485;
			14052: outdata = 32'd51484;
			14053: outdata = 32'd51483;
			14054: outdata = 32'd51482;
			14055: outdata = 32'd51481;
			14056: outdata = 32'd51480;
			14057: outdata = 32'd51479;
			14058: outdata = 32'd51478;
			14059: outdata = 32'd51477;
			14060: outdata = 32'd51476;
			14061: outdata = 32'd51475;
			14062: outdata = 32'd51474;
			14063: outdata = 32'd51473;
			14064: outdata = 32'd51472;
			14065: outdata = 32'd51471;
			14066: outdata = 32'd51470;
			14067: outdata = 32'd51469;
			14068: outdata = 32'd51468;
			14069: outdata = 32'd51467;
			14070: outdata = 32'd51466;
			14071: outdata = 32'd51465;
			14072: outdata = 32'd51464;
			14073: outdata = 32'd51463;
			14074: outdata = 32'd51462;
			14075: outdata = 32'd51461;
			14076: outdata = 32'd51460;
			14077: outdata = 32'd51459;
			14078: outdata = 32'd51458;
			14079: outdata = 32'd51457;
			14080: outdata = 32'd51456;
			14081: outdata = 32'd51455;
			14082: outdata = 32'd51454;
			14083: outdata = 32'd51453;
			14084: outdata = 32'd51452;
			14085: outdata = 32'd51451;
			14086: outdata = 32'd51450;
			14087: outdata = 32'd51449;
			14088: outdata = 32'd51448;
			14089: outdata = 32'd51447;
			14090: outdata = 32'd51446;
			14091: outdata = 32'd51445;
			14092: outdata = 32'd51444;
			14093: outdata = 32'd51443;
			14094: outdata = 32'd51442;
			14095: outdata = 32'd51441;
			14096: outdata = 32'd51440;
			14097: outdata = 32'd51439;
			14098: outdata = 32'd51438;
			14099: outdata = 32'd51437;
			14100: outdata = 32'd51436;
			14101: outdata = 32'd51435;
			14102: outdata = 32'd51434;
			14103: outdata = 32'd51433;
			14104: outdata = 32'd51432;
			14105: outdata = 32'd51431;
			14106: outdata = 32'd51430;
			14107: outdata = 32'd51429;
			14108: outdata = 32'd51428;
			14109: outdata = 32'd51427;
			14110: outdata = 32'd51426;
			14111: outdata = 32'd51425;
			14112: outdata = 32'd51424;
			14113: outdata = 32'd51423;
			14114: outdata = 32'd51422;
			14115: outdata = 32'd51421;
			14116: outdata = 32'd51420;
			14117: outdata = 32'd51419;
			14118: outdata = 32'd51418;
			14119: outdata = 32'd51417;
			14120: outdata = 32'd51416;
			14121: outdata = 32'd51415;
			14122: outdata = 32'd51414;
			14123: outdata = 32'd51413;
			14124: outdata = 32'd51412;
			14125: outdata = 32'd51411;
			14126: outdata = 32'd51410;
			14127: outdata = 32'd51409;
			14128: outdata = 32'd51408;
			14129: outdata = 32'd51407;
			14130: outdata = 32'd51406;
			14131: outdata = 32'd51405;
			14132: outdata = 32'd51404;
			14133: outdata = 32'd51403;
			14134: outdata = 32'd51402;
			14135: outdata = 32'd51401;
			14136: outdata = 32'd51400;
			14137: outdata = 32'd51399;
			14138: outdata = 32'd51398;
			14139: outdata = 32'd51397;
			14140: outdata = 32'd51396;
			14141: outdata = 32'd51395;
			14142: outdata = 32'd51394;
			14143: outdata = 32'd51393;
			14144: outdata = 32'd51392;
			14145: outdata = 32'd51391;
			14146: outdata = 32'd51390;
			14147: outdata = 32'd51389;
			14148: outdata = 32'd51388;
			14149: outdata = 32'd51387;
			14150: outdata = 32'd51386;
			14151: outdata = 32'd51385;
			14152: outdata = 32'd51384;
			14153: outdata = 32'd51383;
			14154: outdata = 32'd51382;
			14155: outdata = 32'd51381;
			14156: outdata = 32'd51380;
			14157: outdata = 32'd51379;
			14158: outdata = 32'd51378;
			14159: outdata = 32'd51377;
			14160: outdata = 32'd51376;
			14161: outdata = 32'd51375;
			14162: outdata = 32'd51374;
			14163: outdata = 32'd51373;
			14164: outdata = 32'd51372;
			14165: outdata = 32'd51371;
			14166: outdata = 32'd51370;
			14167: outdata = 32'd51369;
			14168: outdata = 32'd51368;
			14169: outdata = 32'd51367;
			14170: outdata = 32'd51366;
			14171: outdata = 32'd51365;
			14172: outdata = 32'd51364;
			14173: outdata = 32'd51363;
			14174: outdata = 32'd51362;
			14175: outdata = 32'd51361;
			14176: outdata = 32'd51360;
			14177: outdata = 32'd51359;
			14178: outdata = 32'd51358;
			14179: outdata = 32'd51357;
			14180: outdata = 32'd51356;
			14181: outdata = 32'd51355;
			14182: outdata = 32'd51354;
			14183: outdata = 32'd51353;
			14184: outdata = 32'd51352;
			14185: outdata = 32'd51351;
			14186: outdata = 32'd51350;
			14187: outdata = 32'd51349;
			14188: outdata = 32'd51348;
			14189: outdata = 32'd51347;
			14190: outdata = 32'd51346;
			14191: outdata = 32'd51345;
			14192: outdata = 32'd51344;
			14193: outdata = 32'd51343;
			14194: outdata = 32'd51342;
			14195: outdata = 32'd51341;
			14196: outdata = 32'd51340;
			14197: outdata = 32'd51339;
			14198: outdata = 32'd51338;
			14199: outdata = 32'd51337;
			14200: outdata = 32'd51336;
			14201: outdata = 32'd51335;
			14202: outdata = 32'd51334;
			14203: outdata = 32'd51333;
			14204: outdata = 32'd51332;
			14205: outdata = 32'd51331;
			14206: outdata = 32'd51330;
			14207: outdata = 32'd51329;
			14208: outdata = 32'd51328;
			14209: outdata = 32'd51327;
			14210: outdata = 32'd51326;
			14211: outdata = 32'd51325;
			14212: outdata = 32'd51324;
			14213: outdata = 32'd51323;
			14214: outdata = 32'd51322;
			14215: outdata = 32'd51321;
			14216: outdata = 32'd51320;
			14217: outdata = 32'd51319;
			14218: outdata = 32'd51318;
			14219: outdata = 32'd51317;
			14220: outdata = 32'd51316;
			14221: outdata = 32'd51315;
			14222: outdata = 32'd51314;
			14223: outdata = 32'd51313;
			14224: outdata = 32'd51312;
			14225: outdata = 32'd51311;
			14226: outdata = 32'd51310;
			14227: outdata = 32'd51309;
			14228: outdata = 32'd51308;
			14229: outdata = 32'd51307;
			14230: outdata = 32'd51306;
			14231: outdata = 32'd51305;
			14232: outdata = 32'd51304;
			14233: outdata = 32'd51303;
			14234: outdata = 32'd51302;
			14235: outdata = 32'd51301;
			14236: outdata = 32'd51300;
			14237: outdata = 32'd51299;
			14238: outdata = 32'd51298;
			14239: outdata = 32'd51297;
			14240: outdata = 32'd51296;
			14241: outdata = 32'd51295;
			14242: outdata = 32'd51294;
			14243: outdata = 32'd51293;
			14244: outdata = 32'd51292;
			14245: outdata = 32'd51291;
			14246: outdata = 32'd51290;
			14247: outdata = 32'd51289;
			14248: outdata = 32'd51288;
			14249: outdata = 32'd51287;
			14250: outdata = 32'd51286;
			14251: outdata = 32'd51285;
			14252: outdata = 32'd51284;
			14253: outdata = 32'd51283;
			14254: outdata = 32'd51282;
			14255: outdata = 32'd51281;
			14256: outdata = 32'd51280;
			14257: outdata = 32'd51279;
			14258: outdata = 32'd51278;
			14259: outdata = 32'd51277;
			14260: outdata = 32'd51276;
			14261: outdata = 32'd51275;
			14262: outdata = 32'd51274;
			14263: outdata = 32'd51273;
			14264: outdata = 32'd51272;
			14265: outdata = 32'd51271;
			14266: outdata = 32'd51270;
			14267: outdata = 32'd51269;
			14268: outdata = 32'd51268;
			14269: outdata = 32'd51267;
			14270: outdata = 32'd51266;
			14271: outdata = 32'd51265;
			14272: outdata = 32'd51264;
			14273: outdata = 32'd51263;
			14274: outdata = 32'd51262;
			14275: outdata = 32'd51261;
			14276: outdata = 32'd51260;
			14277: outdata = 32'd51259;
			14278: outdata = 32'd51258;
			14279: outdata = 32'd51257;
			14280: outdata = 32'd51256;
			14281: outdata = 32'd51255;
			14282: outdata = 32'd51254;
			14283: outdata = 32'd51253;
			14284: outdata = 32'd51252;
			14285: outdata = 32'd51251;
			14286: outdata = 32'd51250;
			14287: outdata = 32'd51249;
			14288: outdata = 32'd51248;
			14289: outdata = 32'd51247;
			14290: outdata = 32'd51246;
			14291: outdata = 32'd51245;
			14292: outdata = 32'd51244;
			14293: outdata = 32'd51243;
			14294: outdata = 32'd51242;
			14295: outdata = 32'd51241;
			14296: outdata = 32'd51240;
			14297: outdata = 32'd51239;
			14298: outdata = 32'd51238;
			14299: outdata = 32'd51237;
			14300: outdata = 32'd51236;
			14301: outdata = 32'd51235;
			14302: outdata = 32'd51234;
			14303: outdata = 32'd51233;
			14304: outdata = 32'd51232;
			14305: outdata = 32'd51231;
			14306: outdata = 32'd51230;
			14307: outdata = 32'd51229;
			14308: outdata = 32'd51228;
			14309: outdata = 32'd51227;
			14310: outdata = 32'd51226;
			14311: outdata = 32'd51225;
			14312: outdata = 32'd51224;
			14313: outdata = 32'd51223;
			14314: outdata = 32'd51222;
			14315: outdata = 32'd51221;
			14316: outdata = 32'd51220;
			14317: outdata = 32'd51219;
			14318: outdata = 32'd51218;
			14319: outdata = 32'd51217;
			14320: outdata = 32'd51216;
			14321: outdata = 32'd51215;
			14322: outdata = 32'd51214;
			14323: outdata = 32'd51213;
			14324: outdata = 32'd51212;
			14325: outdata = 32'd51211;
			14326: outdata = 32'd51210;
			14327: outdata = 32'd51209;
			14328: outdata = 32'd51208;
			14329: outdata = 32'd51207;
			14330: outdata = 32'd51206;
			14331: outdata = 32'd51205;
			14332: outdata = 32'd51204;
			14333: outdata = 32'd51203;
			14334: outdata = 32'd51202;
			14335: outdata = 32'd51201;
			14336: outdata = 32'd51200;
			14337: outdata = 32'd51199;
			14338: outdata = 32'd51198;
			14339: outdata = 32'd51197;
			14340: outdata = 32'd51196;
			14341: outdata = 32'd51195;
			14342: outdata = 32'd51194;
			14343: outdata = 32'd51193;
			14344: outdata = 32'd51192;
			14345: outdata = 32'd51191;
			14346: outdata = 32'd51190;
			14347: outdata = 32'd51189;
			14348: outdata = 32'd51188;
			14349: outdata = 32'd51187;
			14350: outdata = 32'd51186;
			14351: outdata = 32'd51185;
			14352: outdata = 32'd51184;
			14353: outdata = 32'd51183;
			14354: outdata = 32'd51182;
			14355: outdata = 32'd51181;
			14356: outdata = 32'd51180;
			14357: outdata = 32'd51179;
			14358: outdata = 32'd51178;
			14359: outdata = 32'd51177;
			14360: outdata = 32'd51176;
			14361: outdata = 32'd51175;
			14362: outdata = 32'd51174;
			14363: outdata = 32'd51173;
			14364: outdata = 32'd51172;
			14365: outdata = 32'd51171;
			14366: outdata = 32'd51170;
			14367: outdata = 32'd51169;
			14368: outdata = 32'd51168;
			14369: outdata = 32'd51167;
			14370: outdata = 32'd51166;
			14371: outdata = 32'd51165;
			14372: outdata = 32'd51164;
			14373: outdata = 32'd51163;
			14374: outdata = 32'd51162;
			14375: outdata = 32'd51161;
			14376: outdata = 32'd51160;
			14377: outdata = 32'd51159;
			14378: outdata = 32'd51158;
			14379: outdata = 32'd51157;
			14380: outdata = 32'd51156;
			14381: outdata = 32'd51155;
			14382: outdata = 32'd51154;
			14383: outdata = 32'd51153;
			14384: outdata = 32'd51152;
			14385: outdata = 32'd51151;
			14386: outdata = 32'd51150;
			14387: outdata = 32'd51149;
			14388: outdata = 32'd51148;
			14389: outdata = 32'd51147;
			14390: outdata = 32'd51146;
			14391: outdata = 32'd51145;
			14392: outdata = 32'd51144;
			14393: outdata = 32'd51143;
			14394: outdata = 32'd51142;
			14395: outdata = 32'd51141;
			14396: outdata = 32'd51140;
			14397: outdata = 32'd51139;
			14398: outdata = 32'd51138;
			14399: outdata = 32'd51137;
			14400: outdata = 32'd51136;
			14401: outdata = 32'd51135;
			14402: outdata = 32'd51134;
			14403: outdata = 32'd51133;
			14404: outdata = 32'd51132;
			14405: outdata = 32'd51131;
			14406: outdata = 32'd51130;
			14407: outdata = 32'd51129;
			14408: outdata = 32'd51128;
			14409: outdata = 32'd51127;
			14410: outdata = 32'd51126;
			14411: outdata = 32'd51125;
			14412: outdata = 32'd51124;
			14413: outdata = 32'd51123;
			14414: outdata = 32'd51122;
			14415: outdata = 32'd51121;
			14416: outdata = 32'd51120;
			14417: outdata = 32'd51119;
			14418: outdata = 32'd51118;
			14419: outdata = 32'd51117;
			14420: outdata = 32'd51116;
			14421: outdata = 32'd51115;
			14422: outdata = 32'd51114;
			14423: outdata = 32'd51113;
			14424: outdata = 32'd51112;
			14425: outdata = 32'd51111;
			14426: outdata = 32'd51110;
			14427: outdata = 32'd51109;
			14428: outdata = 32'd51108;
			14429: outdata = 32'd51107;
			14430: outdata = 32'd51106;
			14431: outdata = 32'd51105;
			14432: outdata = 32'd51104;
			14433: outdata = 32'd51103;
			14434: outdata = 32'd51102;
			14435: outdata = 32'd51101;
			14436: outdata = 32'd51100;
			14437: outdata = 32'd51099;
			14438: outdata = 32'd51098;
			14439: outdata = 32'd51097;
			14440: outdata = 32'd51096;
			14441: outdata = 32'd51095;
			14442: outdata = 32'd51094;
			14443: outdata = 32'd51093;
			14444: outdata = 32'd51092;
			14445: outdata = 32'd51091;
			14446: outdata = 32'd51090;
			14447: outdata = 32'd51089;
			14448: outdata = 32'd51088;
			14449: outdata = 32'd51087;
			14450: outdata = 32'd51086;
			14451: outdata = 32'd51085;
			14452: outdata = 32'd51084;
			14453: outdata = 32'd51083;
			14454: outdata = 32'd51082;
			14455: outdata = 32'd51081;
			14456: outdata = 32'd51080;
			14457: outdata = 32'd51079;
			14458: outdata = 32'd51078;
			14459: outdata = 32'd51077;
			14460: outdata = 32'd51076;
			14461: outdata = 32'd51075;
			14462: outdata = 32'd51074;
			14463: outdata = 32'd51073;
			14464: outdata = 32'd51072;
			14465: outdata = 32'd51071;
			14466: outdata = 32'd51070;
			14467: outdata = 32'd51069;
			14468: outdata = 32'd51068;
			14469: outdata = 32'd51067;
			14470: outdata = 32'd51066;
			14471: outdata = 32'd51065;
			14472: outdata = 32'd51064;
			14473: outdata = 32'd51063;
			14474: outdata = 32'd51062;
			14475: outdata = 32'd51061;
			14476: outdata = 32'd51060;
			14477: outdata = 32'd51059;
			14478: outdata = 32'd51058;
			14479: outdata = 32'd51057;
			14480: outdata = 32'd51056;
			14481: outdata = 32'd51055;
			14482: outdata = 32'd51054;
			14483: outdata = 32'd51053;
			14484: outdata = 32'd51052;
			14485: outdata = 32'd51051;
			14486: outdata = 32'd51050;
			14487: outdata = 32'd51049;
			14488: outdata = 32'd51048;
			14489: outdata = 32'd51047;
			14490: outdata = 32'd51046;
			14491: outdata = 32'd51045;
			14492: outdata = 32'd51044;
			14493: outdata = 32'd51043;
			14494: outdata = 32'd51042;
			14495: outdata = 32'd51041;
			14496: outdata = 32'd51040;
			14497: outdata = 32'd51039;
			14498: outdata = 32'd51038;
			14499: outdata = 32'd51037;
			14500: outdata = 32'd51036;
			14501: outdata = 32'd51035;
			14502: outdata = 32'd51034;
			14503: outdata = 32'd51033;
			14504: outdata = 32'd51032;
			14505: outdata = 32'd51031;
			14506: outdata = 32'd51030;
			14507: outdata = 32'd51029;
			14508: outdata = 32'd51028;
			14509: outdata = 32'd51027;
			14510: outdata = 32'd51026;
			14511: outdata = 32'd51025;
			14512: outdata = 32'd51024;
			14513: outdata = 32'd51023;
			14514: outdata = 32'd51022;
			14515: outdata = 32'd51021;
			14516: outdata = 32'd51020;
			14517: outdata = 32'd51019;
			14518: outdata = 32'd51018;
			14519: outdata = 32'd51017;
			14520: outdata = 32'd51016;
			14521: outdata = 32'd51015;
			14522: outdata = 32'd51014;
			14523: outdata = 32'd51013;
			14524: outdata = 32'd51012;
			14525: outdata = 32'd51011;
			14526: outdata = 32'd51010;
			14527: outdata = 32'd51009;
			14528: outdata = 32'd51008;
			14529: outdata = 32'd51007;
			14530: outdata = 32'd51006;
			14531: outdata = 32'd51005;
			14532: outdata = 32'd51004;
			14533: outdata = 32'd51003;
			14534: outdata = 32'd51002;
			14535: outdata = 32'd51001;
			14536: outdata = 32'd51000;
			14537: outdata = 32'd50999;
			14538: outdata = 32'd50998;
			14539: outdata = 32'd50997;
			14540: outdata = 32'd50996;
			14541: outdata = 32'd50995;
			14542: outdata = 32'd50994;
			14543: outdata = 32'd50993;
			14544: outdata = 32'd50992;
			14545: outdata = 32'd50991;
			14546: outdata = 32'd50990;
			14547: outdata = 32'd50989;
			14548: outdata = 32'd50988;
			14549: outdata = 32'd50987;
			14550: outdata = 32'd50986;
			14551: outdata = 32'd50985;
			14552: outdata = 32'd50984;
			14553: outdata = 32'd50983;
			14554: outdata = 32'd50982;
			14555: outdata = 32'd50981;
			14556: outdata = 32'd50980;
			14557: outdata = 32'd50979;
			14558: outdata = 32'd50978;
			14559: outdata = 32'd50977;
			14560: outdata = 32'd50976;
			14561: outdata = 32'd50975;
			14562: outdata = 32'd50974;
			14563: outdata = 32'd50973;
			14564: outdata = 32'd50972;
			14565: outdata = 32'd50971;
			14566: outdata = 32'd50970;
			14567: outdata = 32'd50969;
			14568: outdata = 32'd50968;
			14569: outdata = 32'd50967;
			14570: outdata = 32'd50966;
			14571: outdata = 32'd50965;
			14572: outdata = 32'd50964;
			14573: outdata = 32'd50963;
			14574: outdata = 32'd50962;
			14575: outdata = 32'd50961;
			14576: outdata = 32'd50960;
			14577: outdata = 32'd50959;
			14578: outdata = 32'd50958;
			14579: outdata = 32'd50957;
			14580: outdata = 32'd50956;
			14581: outdata = 32'd50955;
			14582: outdata = 32'd50954;
			14583: outdata = 32'd50953;
			14584: outdata = 32'd50952;
			14585: outdata = 32'd50951;
			14586: outdata = 32'd50950;
			14587: outdata = 32'd50949;
			14588: outdata = 32'd50948;
			14589: outdata = 32'd50947;
			14590: outdata = 32'd50946;
			14591: outdata = 32'd50945;
			14592: outdata = 32'd50944;
			14593: outdata = 32'd50943;
			14594: outdata = 32'd50942;
			14595: outdata = 32'd50941;
			14596: outdata = 32'd50940;
			14597: outdata = 32'd50939;
			14598: outdata = 32'd50938;
			14599: outdata = 32'd50937;
			14600: outdata = 32'd50936;
			14601: outdata = 32'd50935;
			14602: outdata = 32'd50934;
			14603: outdata = 32'd50933;
			14604: outdata = 32'd50932;
			14605: outdata = 32'd50931;
			14606: outdata = 32'd50930;
			14607: outdata = 32'd50929;
			14608: outdata = 32'd50928;
			14609: outdata = 32'd50927;
			14610: outdata = 32'd50926;
			14611: outdata = 32'd50925;
			14612: outdata = 32'd50924;
			14613: outdata = 32'd50923;
			14614: outdata = 32'd50922;
			14615: outdata = 32'd50921;
			14616: outdata = 32'd50920;
			14617: outdata = 32'd50919;
			14618: outdata = 32'd50918;
			14619: outdata = 32'd50917;
			14620: outdata = 32'd50916;
			14621: outdata = 32'd50915;
			14622: outdata = 32'd50914;
			14623: outdata = 32'd50913;
			14624: outdata = 32'd50912;
			14625: outdata = 32'd50911;
			14626: outdata = 32'd50910;
			14627: outdata = 32'd50909;
			14628: outdata = 32'd50908;
			14629: outdata = 32'd50907;
			14630: outdata = 32'd50906;
			14631: outdata = 32'd50905;
			14632: outdata = 32'd50904;
			14633: outdata = 32'd50903;
			14634: outdata = 32'd50902;
			14635: outdata = 32'd50901;
			14636: outdata = 32'd50900;
			14637: outdata = 32'd50899;
			14638: outdata = 32'd50898;
			14639: outdata = 32'd50897;
			14640: outdata = 32'd50896;
			14641: outdata = 32'd50895;
			14642: outdata = 32'd50894;
			14643: outdata = 32'd50893;
			14644: outdata = 32'd50892;
			14645: outdata = 32'd50891;
			14646: outdata = 32'd50890;
			14647: outdata = 32'd50889;
			14648: outdata = 32'd50888;
			14649: outdata = 32'd50887;
			14650: outdata = 32'd50886;
			14651: outdata = 32'd50885;
			14652: outdata = 32'd50884;
			14653: outdata = 32'd50883;
			14654: outdata = 32'd50882;
			14655: outdata = 32'd50881;
			14656: outdata = 32'd50880;
			14657: outdata = 32'd50879;
			14658: outdata = 32'd50878;
			14659: outdata = 32'd50877;
			14660: outdata = 32'd50876;
			14661: outdata = 32'd50875;
			14662: outdata = 32'd50874;
			14663: outdata = 32'd50873;
			14664: outdata = 32'd50872;
			14665: outdata = 32'd50871;
			14666: outdata = 32'd50870;
			14667: outdata = 32'd50869;
			14668: outdata = 32'd50868;
			14669: outdata = 32'd50867;
			14670: outdata = 32'd50866;
			14671: outdata = 32'd50865;
			14672: outdata = 32'd50864;
			14673: outdata = 32'd50863;
			14674: outdata = 32'd50862;
			14675: outdata = 32'd50861;
			14676: outdata = 32'd50860;
			14677: outdata = 32'd50859;
			14678: outdata = 32'd50858;
			14679: outdata = 32'd50857;
			14680: outdata = 32'd50856;
			14681: outdata = 32'd50855;
			14682: outdata = 32'd50854;
			14683: outdata = 32'd50853;
			14684: outdata = 32'd50852;
			14685: outdata = 32'd50851;
			14686: outdata = 32'd50850;
			14687: outdata = 32'd50849;
			14688: outdata = 32'd50848;
			14689: outdata = 32'd50847;
			14690: outdata = 32'd50846;
			14691: outdata = 32'd50845;
			14692: outdata = 32'd50844;
			14693: outdata = 32'd50843;
			14694: outdata = 32'd50842;
			14695: outdata = 32'd50841;
			14696: outdata = 32'd50840;
			14697: outdata = 32'd50839;
			14698: outdata = 32'd50838;
			14699: outdata = 32'd50837;
			14700: outdata = 32'd50836;
			14701: outdata = 32'd50835;
			14702: outdata = 32'd50834;
			14703: outdata = 32'd50833;
			14704: outdata = 32'd50832;
			14705: outdata = 32'd50831;
			14706: outdata = 32'd50830;
			14707: outdata = 32'd50829;
			14708: outdata = 32'd50828;
			14709: outdata = 32'd50827;
			14710: outdata = 32'd50826;
			14711: outdata = 32'd50825;
			14712: outdata = 32'd50824;
			14713: outdata = 32'd50823;
			14714: outdata = 32'd50822;
			14715: outdata = 32'd50821;
			14716: outdata = 32'd50820;
			14717: outdata = 32'd50819;
			14718: outdata = 32'd50818;
			14719: outdata = 32'd50817;
			14720: outdata = 32'd50816;
			14721: outdata = 32'd50815;
			14722: outdata = 32'd50814;
			14723: outdata = 32'd50813;
			14724: outdata = 32'd50812;
			14725: outdata = 32'd50811;
			14726: outdata = 32'd50810;
			14727: outdata = 32'd50809;
			14728: outdata = 32'd50808;
			14729: outdata = 32'd50807;
			14730: outdata = 32'd50806;
			14731: outdata = 32'd50805;
			14732: outdata = 32'd50804;
			14733: outdata = 32'd50803;
			14734: outdata = 32'd50802;
			14735: outdata = 32'd50801;
			14736: outdata = 32'd50800;
			14737: outdata = 32'd50799;
			14738: outdata = 32'd50798;
			14739: outdata = 32'd50797;
			14740: outdata = 32'd50796;
			14741: outdata = 32'd50795;
			14742: outdata = 32'd50794;
			14743: outdata = 32'd50793;
			14744: outdata = 32'd50792;
			14745: outdata = 32'd50791;
			14746: outdata = 32'd50790;
			14747: outdata = 32'd50789;
			14748: outdata = 32'd50788;
			14749: outdata = 32'd50787;
			14750: outdata = 32'd50786;
			14751: outdata = 32'd50785;
			14752: outdata = 32'd50784;
			14753: outdata = 32'd50783;
			14754: outdata = 32'd50782;
			14755: outdata = 32'd50781;
			14756: outdata = 32'd50780;
			14757: outdata = 32'd50779;
			14758: outdata = 32'd50778;
			14759: outdata = 32'd50777;
			14760: outdata = 32'd50776;
			14761: outdata = 32'd50775;
			14762: outdata = 32'd50774;
			14763: outdata = 32'd50773;
			14764: outdata = 32'd50772;
			14765: outdata = 32'd50771;
			14766: outdata = 32'd50770;
			14767: outdata = 32'd50769;
			14768: outdata = 32'd50768;
			14769: outdata = 32'd50767;
			14770: outdata = 32'd50766;
			14771: outdata = 32'd50765;
			14772: outdata = 32'd50764;
			14773: outdata = 32'd50763;
			14774: outdata = 32'd50762;
			14775: outdata = 32'd50761;
			14776: outdata = 32'd50760;
			14777: outdata = 32'd50759;
			14778: outdata = 32'd50758;
			14779: outdata = 32'd50757;
			14780: outdata = 32'd50756;
			14781: outdata = 32'd50755;
			14782: outdata = 32'd50754;
			14783: outdata = 32'd50753;
			14784: outdata = 32'd50752;
			14785: outdata = 32'd50751;
			14786: outdata = 32'd50750;
			14787: outdata = 32'd50749;
			14788: outdata = 32'd50748;
			14789: outdata = 32'd50747;
			14790: outdata = 32'd50746;
			14791: outdata = 32'd50745;
			14792: outdata = 32'd50744;
			14793: outdata = 32'd50743;
			14794: outdata = 32'd50742;
			14795: outdata = 32'd50741;
			14796: outdata = 32'd50740;
			14797: outdata = 32'd50739;
			14798: outdata = 32'd50738;
			14799: outdata = 32'd50737;
			14800: outdata = 32'd50736;
			14801: outdata = 32'd50735;
			14802: outdata = 32'd50734;
			14803: outdata = 32'd50733;
			14804: outdata = 32'd50732;
			14805: outdata = 32'd50731;
			14806: outdata = 32'd50730;
			14807: outdata = 32'd50729;
			14808: outdata = 32'd50728;
			14809: outdata = 32'd50727;
			14810: outdata = 32'd50726;
			14811: outdata = 32'd50725;
			14812: outdata = 32'd50724;
			14813: outdata = 32'd50723;
			14814: outdata = 32'd50722;
			14815: outdata = 32'd50721;
			14816: outdata = 32'd50720;
			14817: outdata = 32'd50719;
			14818: outdata = 32'd50718;
			14819: outdata = 32'd50717;
			14820: outdata = 32'd50716;
			14821: outdata = 32'd50715;
			14822: outdata = 32'd50714;
			14823: outdata = 32'd50713;
			14824: outdata = 32'd50712;
			14825: outdata = 32'd50711;
			14826: outdata = 32'd50710;
			14827: outdata = 32'd50709;
			14828: outdata = 32'd50708;
			14829: outdata = 32'd50707;
			14830: outdata = 32'd50706;
			14831: outdata = 32'd50705;
			14832: outdata = 32'd50704;
			14833: outdata = 32'd50703;
			14834: outdata = 32'd50702;
			14835: outdata = 32'd50701;
			14836: outdata = 32'd50700;
			14837: outdata = 32'd50699;
			14838: outdata = 32'd50698;
			14839: outdata = 32'd50697;
			14840: outdata = 32'd50696;
			14841: outdata = 32'd50695;
			14842: outdata = 32'd50694;
			14843: outdata = 32'd50693;
			14844: outdata = 32'd50692;
			14845: outdata = 32'd50691;
			14846: outdata = 32'd50690;
			14847: outdata = 32'd50689;
			14848: outdata = 32'd50688;
			14849: outdata = 32'd50687;
			14850: outdata = 32'd50686;
			14851: outdata = 32'd50685;
			14852: outdata = 32'd50684;
			14853: outdata = 32'd50683;
			14854: outdata = 32'd50682;
			14855: outdata = 32'd50681;
			14856: outdata = 32'd50680;
			14857: outdata = 32'd50679;
			14858: outdata = 32'd50678;
			14859: outdata = 32'd50677;
			14860: outdata = 32'd50676;
			14861: outdata = 32'd50675;
			14862: outdata = 32'd50674;
			14863: outdata = 32'd50673;
			14864: outdata = 32'd50672;
			14865: outdata = 32'd50671;
			14866: outdata = 32'd50670;
			14867: outdata = 32'd50669;
			14868: outdata = 32'd50668;
			14869: outdata = 32'd50667;
			14870: outdata = 32'd50666;
			14871: outdata = 32'd50665;
			14872: outdata = 32'd50664;
			14873: outdata = 32'd50663;
			14874: outdata = 32'd50662;
			14875: outdata = 32'd50661;
			14876: outdata = 32'd50660;
			14877: outdata = 32'd50659;
			14878: outdata = 32'd50658;
			14879: outdata = 32'd50657;
			14880: outdata = 32'd50656;
			14881: outdata = 32'd50655;
			14882: outdata = 32'd50654;
			14883: outdata = 32'd50653;
			14884: outdata = 32'd50652;
			14885: outdata = 32'd50651;
			14886: outdata = 32'd50650;
			14887: outdata = 32'd50649;
			14888: outdata = 32'd50648;
			14889: outdata = 32'd50647;
			14890: outdata = 32'd50646;
			14891: outdata = 32'd50645;
			14892: outdata = 32'd50644;
			14893: outdata = 32'd50643;
			14894: outdata = 32'd50642;
			14895: outdata = 32'd50641;
			14896: outdata = 32'd50640;
			14897: outdata = 32'd50639;
			14898: outdata = 32'd50638;
			14899: outdata = 32'd50637;
			14900: outdata = 32'd50636;
			14901: outdata = 32'd50635;
			14902: outdata = 32'd50634;
			14903: outdata = 32'd50633;
			14904: outdata = 32'd50632;
			14905: outdata = 32'd50631;
			14906: outdata = 32'd50630;
			14907: outdata = 32'd50629;
			14908: outdata = 32'd50628;
			14909: outdata = 32'd50627;
			14910: outdata = 32'd50626;
			14911: outdata = 32'd50625;
			14912: outdata = 32'd50624;
			14913: outdata = 32'd50623;
			14914: outdata = 32'd50622;
			14915: outdata = 32'd50621;
			14916: outdata = 32'd50620;
			14917: outdata = 32'd50619;
			14918: outdata = 32'd50618;
			14919: outdata = 32'd50617;
			14920: outdata = 32'd50616;
			14921: outdata = 32'd50615;
			14922: outdata = 32'd50614;
			14923: outdata = 32'd50613;
			14924: outdata = 32'd50612;
			14925: outdata = 32'd50611;
			14926: outdata = 32'd50610;
			14927: outdata = 32'd50609;
			14928: outdata = 32'd50608;
			14929: outdata = 32'd50607;
			14930: outdata = 32'd50606;
			14931: outdata = 32'd50605;
			14932: outdata = 32'd50604;
			14933: outdata = 32'd50603;
			14934: outdata = 32'd50602;
			14935: outdata = 32'd50601;
			14936: outdata = 32'd50600;
			14937: outdata = 32'd50599;
			14938: outdata = 32'd50598;
			14939: outdata = 32'd50597;
			14940: outdata = 32'd50596;
			14941: outdata = 32'd50595;
			14942: outdata = 32'd50594;
			14943: outdata = 32'd50593;
			14944: outdata = 32'd50592;
			14945: outdata = 32'd50591;
			14946: outdata = 32'd50590;
			14947: outdata = 32'd50589;
			14948: outdata = 32'd50588;
			14949: outdata = 32'd50587;
			14950: outdata = 32'd50586;
			14951: outdata = 32'd50585;
			14952: outdata = 32'd50584;
			14953: outdata = 32'd50583;
			14954: outdata = 32'd50582;
			14955: outdata = 32'd50581;
			14956: outdata = 32'd50580;
			14957: outdata = 32'd50579;
			14958: outdata = 32'd50578;
			14959: outdata = 32'd50577;
			14960: outdata = 32'd50576;
			14961: outdata = 32'd50575;
			14962: outdata = 32'd50574;
			14963: outdata = 32'd50573;
			14964: outdata = 32'd50572;
			14965: outdata = 32'd50571;
			14966: outdata = 32'd50570;
			14967: outdata = 32'd50569;
			14968: outdata = 32'd50568;
			14969: outdata = 32'd50567;
			14970: outdata = 32'd50566;
			14971: outdata = 32'd50565;
			14972: outdata = 32'd50564;
			14973: outdata = 32'd50563;
			14974: outdata = 32'd50562;
			14975: outdata = 32'd50561;
			14976: outdata = 32'd50560;
			14977: outdata = 32'd50559;
			14978: outdata = 32'd50558;
			14979: outdata = 32'd50557;
			14980: outdata = 32'd50556;
			14981: outdata = 32'd50555;
			14982: outdata = 32'd50554;
			14983: outdata = 32'd50553;
			14984: outdata = 32'd50552;
			14985: outdata = 32'd50551;
			14986: outdata = 32'd50550;
			14987: outdata = 32'd50549;
			14988: outdata = 32'd50548;
			14989: outdata = 32'd50547;
			14990: outdata = 32'd50546;
			14991: outdata = 32'd50545;
			14992: outdata = 32'd50544;
			14993: outdata = 32'd50543;
			14994: outdata = 32'd50542;
			14995: outdata = 32'd50541;
			14996: outdata = 32'd50540;
			14997: outdata = 32'd50539;
			14998: outdata = 32'd50538;
			14999: outdata = 32'd50537;
			15000: outdata = 32'd50536;
			15001: outdata = 32'd50535;
			15002: outdata = 32'd50534;
			15003: outdata = 32'd50533;
			15004: outdata = 32'd50532;
			15005: outdata = 32'd50531;
			15006: outdata = 32'd50530;
			15007: outdata = 32'd50529;
			15008: outdata = 32'd50528;
			15009: outdata = 32'd50527;
			15010: outdata = 32'd50526;
			15011: outdata = 32'd50525;
			15012: outdata = 32'd50524;
			15013: outdata = 32'd50523;
			15014: outdata = 32'd50522;
			15015: outdata = 32'd50521;
			15016: outdata = 32'd50520;
			15017: outdata = 32'd50519;
			15018: outdata = 32'd50518;
			15019: outdata = 32'd50517;
			15020: outdata = 32'd50516;
			15021: outdata = 32'd50515;
			15022: outdata = 32'd50514;
			15023: outdata = 32'd50513;
			15024: outdata = 32'd50512;
			15025: outdata = 32'd50511;
			15026: outdata = 32'd50510;
			15027: outdata = 32'd50509;
			15028: outdata = 32'd50508;
			15029: outdata = 32'd50507;
			15030: outdata = 32'd50506;
			15031: outdata = 32'd50505;
			15032: outdata = 32'd50504;
			15033: outdata = 32'd50503;
			15034: outdata = 32'd50502;
			15035: outdata = 32'd50501;
			15036: outdata = 32'd50500;
			15037: outdata = 32'd50499;
			15038: outdata = 32'd50498;
			15039: outdata = 32'd50497;
			15040: outdata = 32'd50496;
			15041: outdata = 32'd50495;
			15042: outdata = 32'd50494;
			15043: outdata = 32'd50493;
			15044: outdata = 32'd50492;
			15045: outdata = 32'd50491;
			15046: outdata = 32'd50490;
			15047: outdata = 32'd50489;
			15048: outdata = 32'd50488;
			15049: outdata = 32'd50487;
			15050: outdata = 32'd50486;
			15051: outdata = 32'd50485;
			15052: outdata = 32'd50484;
			15053: outdata = 32'd50483;
			15054: outdata = 32'd50482;
			15055: outdata = 32'd50481;
			15056: outdata = 32'd50480;
			15057: outdata = 32'd50479;
			15058: outdata = 32'd50478;
			15059: outdata = 32'd50477;
			15060: outdata = 32'd50476;
			15061: outdata = 32'd50475;
			15062: outdata = 32'd50474;
			15063: outdata = 32'd50473;
			15064: outdata = 32'd50472;
			15065: outdata = 32'd50471;
			15066: outdata = 32'd50470;
			15067: outdata = 32'd50469;
			15068: outdata = 32'd50468;
			15069: outdata = 32'd50467;
			15070: outdata = 32'd50466;
			15071: outdata = 32'd50465;
			15072: outdata = 32'd50464;
			15073: outdata = 32'd50463;
			15074: outdata = 32'd50462;
			15075: outdata = 32'd50461;
			15076: outdata = 32'd50460;
			15077: outdata = 32'd50459;
			15078: outdata = 32'd50458;
			15079: outdata = 32'd50457;
			15080: outdata = 32'd50456;
			15081: outdata = 32'd50455;
			15082: outdata = 32'd50454;
			15083: outdata = 32'd50453;
			15084: outdata = 32'd50452;
			15085: outdata = 32'd50451;
			15086: outdata = 32'd50450;
			15087: outdata = 32'd50449;
			15088: outdata = 32'd50448;
			15089: outdata = 32'd50447;
			15090: outdata = 32'd50446;
			15091: outdata = 32'd50445;
			15092: outdata = 32'd50444;
			15093: outdata = 32'd50443;
			15094: outdata = 32'd50442;
			15095: outdata = 32'd50441;
			15096: outdata = 32'd50440;
			15097: outdata = 32'd50439;
			15098: outdata = 32'd50438;
			15099: outdata = 32'd50437;
			15100: outdata = 32'd50436;
			15101: outdata = 32'd50435;
			15102: outdata = 32'd50434;
			15103: outdata = 32'd50433;
			15104: outdata = 32'd50432;
			15105: outdata = 32'd50431;
			15106: outdata = 32'd50430;
			15107: outdata = 32'd50429;
			15108: outdata = 32'd50428;
			15109: outdata = 32'd50427;
			15110: outdata = 32'd50426;
			15111: outdata = 32'd50425;
			15112: outdata = 32'd50424;
			15113: outdata = 32'd50423;
			15114: outdata = 32'd50422;
			15115: outdata = 32'd50421;
			15116: outdata = 32'd50420;
			15117: outdata = 32'd50419;
			15118: outdata = 32'd50418;
			15119: outdata = 32'd50417;
			15120: outdata = 32'd50416;
			15121: outdata = 32'd50415;
			15122: outdata = 32'd50414;
			15123: outdata = 32'd50413;
			15124: outdata = 32'd50412;
			15125: outdata = 32'd50411;
			15126: outdata = 32'd50410;
			15127: outdata = 32'd50409;
			15128: outdata = 32'd50408;
			15129: outdata = 32'd50407;
			15130: outdata = 32'd50406;
			15131: outdata = 32'd50405;
			15132: outdata = 32'd50404;
			15133: outdata = 32'd50403;
			15134: outdata = 32'd50402;
			15135: outdata = 32'd50401;
			15136: outdata = 32'd50400;
			15137: outdata = 32'd50399;
			15138: outdata = 32'd50398;
			15139: outdata = 32'd50397;
			15140: outdata = 32'd50396;
			15141: outdata = 32'd50395;
			15142: outdata = 32'd50394;
			15143: outdata = 32'd50393;
			15144: outdata = 32'd50392;
			15145: outdata = 32'd50391;
			15146: outdata = 32'd50390;
			15147: outdata = 32'd50389;
			15148: outdata = 32'd50388;
			15149: outdata = 32'd50387;
			15150: outdata = 32'd50386;
			15151: outdata = 32'd50385;
			15152: outdata = 32'd50384;
			15153: outdata = 32'd50383;
			15154: outdata = 32'd50382;
			15155: outdata = 32'd50381;
			15156: outdata = 32'd50380;
			15157: outdata = 32'd50379;
			15158: outdata = 32'd50378;
			15159: outdata = 32'd50377;
			15160: outdata = 32'd50376;
			15161: outdata = 32'd50375;
			15162: outdata = 32'd50374;
			15163: outdata = 32'd50373;
			15164: outdata = 32'd50372;
			15165: outdata = 32'd50371;
			15166: outdata = 32'd50370;
			15167: outdata = 32'd50369;
			15168: outdata = 32'd50368;
			15169: outdata = 32'd50367;
			15170: outdata = 32'd50366;
			15171: outdata = 32'd50365;
			15172: outdata = 32'd50364;
			15173: outdata = 32'd50363;
			15174: outdata = 32'd50362;
			15175: outdata = 32'd50361;
			15176: outdata = 32'd50360;
			15177: outdata = 32'd50359;
			15178: outdata = 32'd50358;
			15179: outdata = 32'd50357;
			15180: outdata = 32'd50356;
			15181: outdata = 32'd50355;
			15182: outdata = 32'd50354;
			15183: outdata = 32'd50353;
			15184: outdata = 32'd50352;
			15185: outdata = 32'd50351;
			15186: outdata = 32'd50350;
			15187: outdata = 32'd50349;
			15188: outdata = 32'd50348;
			15189: outdata = 32'd50347;
			15190: outdata = 32'd50346;
			15191: outdata = 32'd50345;
			15192: outdata = 32'd50344;
			15193: outdata = 32'd50343;
			15194: outdata = 32'd50342;
			15195: outdata = 32'd50341;
			15196: outdata = 32'd50340;
			15197: outdata = 32'd50339;
			15198: outdata = 32'd50338;
			15199: outdata = 32'd50337;
			15200: outdata = 32'd50336;
			15201: outdata = 32'd50335;
			15202: outdata = 32'd50334;
			15203: outdata = 32'd50333;
			15204: outdata = 32'd50332;
			15205: outdata = 32'd50331;
			15206: outdata = 32'd50330;
			15207: outdata = 32'd50329;
			15208: outdata = 32'd50328;
			15209: outdata = 32'd50327;
			15210: outdata = 32'd50326;
			15211: outdata = 32'd50325;
			15212: outdata = 32'd50324;
			15213: outdata = 32'd50323;
			15214: outdata = 32'd50322;
			15215: outdata = 32'd50321;
			15216: outdata = 32'd50320;
			15217: outdata = 32'd50319;
			15218: outdata = 32'd50318;
			15219: outdata = 32'd50317;
			15220: outdata = 32'd50316;
			15221: outdata = 32'd50315;
			15222: outdata = 32'd50314;
			15223: outdata = 32'd50313;
			15224: outdata = 32'd50312;
			15225: outdata = 32'd50311;
			15226: outdata = 32'd50310;
			15227: outdata = 32'd50309;
			15228: outdata = 32'd50308;
			15229: outdata = 32'd50307;
			15230: outdata = 32'd50306;
			15231: outdata = 32'd50305;
			15232: outdata = 32'd50304;
			15233: outdata = 32'd50303;
			15234: outdata = 32'd50302;
			15235: outdata = 32'd50301;
			15236: outdata = 32'd50300;
			15237: outdata = 32'd50299;
			15238: outdata = 32'd50298;
			15239: outdata = 32'd50297;
			15240: outdata = 32'd50296;
			15241: outdata = 32'd50295;
			15242: outdata = 32'd50294;
			15243: outdata = 32'd50293;
			15244: outdata = 32'd50292;
			15245: outdata = 32'd50291;
			15246: outdata = 32'd50290;
			15247: outdata = 32'd50289;
			15248: outdata = 32'd50288;
			15249: outdata = 32'd50287;
			15250: outdata = 32'd50286;
			15251: outdata = 32'd50285;
			15252: outdata = 32'd50284;
			15253: outdata = 32'd50283;
			15254: outdata = 32'd50282;
			15255: outdata = 32'd50281;
			15256: outdata = 32'd50280;
			15257: outdata = 32'd50279;
			15258: outdata = 32'd50278;
			15259: outdata = 32'd50277;
			15260: outdata = 32'd50276;
			15261: outdata = 32'd50275;
			15262: outdata = 32'd50274;
			15263: outdata = 32'd50273;
			15264: outdata = 32'd50272;
			15265: outdata = 32'd50271;
			15266: outdata = 32'd50270;
			15267: outdata = 32'd50269;
			15268: outdata = 32'd50268;
			15269: outdata = 32'd50267;
			15270: outdata = 32'd50266;
			15271: outdata = 32'd50265;
			15272: outdata = 32'd50264;
			15273: outdata = 32'd50263;
			15274: outdata = 32'd50262;
			15275: outdata = 32'd50261;
			15276: outdata = 32'd50260;
			15277: outdata = 32'd50259;
			15278: outdata = 32'd50258;
			15279: outdata = 32'd50257;
			15280: outdata = 32'd50256;
			15281: outdata = 32'd50255;
			15282: outdata = 32'd50254;
			15283: outdata = 32'd50253;
			15284: outdata = 32'd50252;
			15285: outdata = 32'd50251;
			15286: outdata = 32'd50250;
			15287: outdata = 32'd50249;
			15288: outdata = 32'd50248;
			15289: outdata = 32'd50247;
			15290: outdata = 32'd50246;
			15291: outdata = 32'd50245;
			15292: outdata = 32'd50244;
			15293: outdata = 32'd50243;
			15294: outdata = 32'd50242;
			15295: outdata = 32'd50241;
			15296: outdata = 32'd50240;
			15297: outdata = 32'd50239;
			15298: outdata = 32'd50238;
			15299: outdata = 32'd50237;
			15300: outdata = 32'd50236;
			15301: outdata = 32'd50235;
			15302: outdata = 32'd50234;
			15303: outdata = 32'd50233;
			15304: outdata = 32'd50232;
			15305: outdata = 32'd50231;
			15306: outdata = 32'd50230;
			15307: outdata = 32'd50229;
			15308: outdata = 32'd50228;
			15309: outdata = 32'd50227;
			15310: outdata = 32'd50226;
			15311: outdata = 32'd50225;
			15312: outdata = 32'd50224;
			15313: outdata = 32'd50223;
			15314: outdata = 32'd50222;
			15315: outdata = 32'd50221;
			15316: outdata = 32'd50220;
			15317: outdata = 32'd50219;
			15318: outdata = 32'd50218;
			15319: outdata = 32'd50217;
			15320: outdata = 32'd50216;
			15321: outdata = 32'd50215;
			15322: outdata = 32'd50214;
			15323: outdata = 32'd50213;
			15324: outdata = 32'd50212;
			15325: outdata = 32'd50211;
			15326: outdata = 32'd50210;
			15327: outdata = 32'd50209;
			15328: outdata = 32'd50208;
			15329: outdata = 32'd50207;
			15330: outdata = 32'd50206;
			15331: outdata = 32'd50205;
			15332: outdata = 32'd50204;
			15333: outdata = 32'd50203;
			15334: outdata = 32'd50202;
			15335: outdata = 32'd50201;
			15336: outdata = 32'd50200;
			15337: outdata = 32'd50199;
			15338: outdata = 32'd50198;
			15339: outdata = 32'd50197;
			15340: outdata = 32'd50196;
			15341: outdata = 32'd50195;
			15342: outdata = 32'd50194;
			15343: outdata = 32'd50193;
			15344: outdata = 32'd50192;
			15345: outdata = 32'd50191;
			15346: outdata = 32'd50190;
			15347: outdata = 32'd50189;
			15348: outdata = 32'd50188;
			15349: outdata = 32'd50187;
			15350: outdata = 32'd50186;
			15351: outdata = 32'd50185;
			15352: outdata = 32'd50184;
			15353: outdata = 32'd50183;
			15354: outdata = 32'd50182;
			15355: outdata = 32'd50181;
			15356: outdata = 32'd50180;
			15357: outdata = 32'd50179;
			15358: outdata = 32'd50178;
			15359: outdata = 32'd50177;
			15360: outdata = 32'd50176;
			15361: outdata = 32'd50175;
			15362: outdata = 32'd50174;
			15363: outdata = 32'd50173;
			15364: outdata = 32'd50172;
			15365: outdata = 32'd50171;
			15366: outdata = 32'd50170;
			15367: outdata = 32'd50169;
			15368: outdata = 32'd50168;
			15369: outdata = 32'd50167;
			15370: outdata = 32'd50166;
			15371: outdata = 32'd50165;
			15372: outdata = 32'd50164;
			15373: outdata = 32'd50163;
			15374: outdata = 32'd50162;
			15375: outdata = 32'd50161;
			15376: outdata = 32'd50160;
			15377: outdata = 32'd50159;
			15378: outdata = 32'd50158;
			15379: outdata = 32'd50157;
			15380: outdata = 32'd50156;
			15381: outdata = 32'd50155;
			15382: outdata = 32'd50154;
			15383: outdata = 32'd50153;
			15384: outdata = 32'd50152;
			15385: outdata = 32'd50151;
			15386: outdata = 32'd50150;
			15387: outdata = 32'd50149;
			15388: outdata = 32'd50148;
			15389: outdata = 32'd50147;
			15390: outdata = 32'd50146;
			15391: outdata = 32'd50145;
			15392: outdata = 32'd50144;
			15393: outdata = 32'd50143;
			15394: outdata = 32'd50142;
			15395: outdata = 32'd50141;
			15396: outdata = 32'd50140;
			15397: outdata = 32'd50139;
			15398: outdata = 32'd50138;
			15399: outdata = 32'd50137;
			15400: outdata = 32'd50136;
			15401: outdata = 32'd50135;
			15402: outdata = 32'd50134;
			15403: outdata = 32'd50133;
			15404: outdata = 32'd50132;
			15405: outdata = 32'd50131;
			15406: outdata = 32'd50130;
			15407: outdata = 32'd50129;
			15408: outdata = 32'd50128;
			15409: outdata = 32'd50127;
			15410: outdata = 32'd50126;
			15411: outdata = 32'd50125;
			15412: outdata = 32'd50124;
			15413: outdata = 32'd50123;
			15414: outdata = 32'd50122;
			15415: outdata = 32'd50121;
			15416: outdata = 32'd50120;
			15417: outdata = 32'd50119;
			15418: outdata = 32'd50118;
			15419: outdata = 32'd50117;
			15420: outdata = 32'd50116;
			15421: outdata = 32'd50115;
			15422: outdata = 32'd50114;
			15423: outdata = 32'd50113;
			15424: outdata = 32'd50112;
			15425: outdata = 32'd50111;
			15426: outdata = 32'd50110;
			15427: outdata = 32'd50109;
			15428: outdata = 32'd50108;
			15429: outdata = 32'd50107;
			15430: outdata = 32'd50106;
			15431: outdata = 32'd50105;
			15432: outdata = 32'd50104;
			15433: outdata = 32'd50103;
			15434: outdata = 32'd50102;
			15435: outdata = 32'd50101;
			15436: outdata = 32'd50100;
			15437: outdata = 32'd50099;
			15438: outdata = 32'd50098;
			15439: outdata = 32'd50097;
			15440: outdata = 32'd50096;
			15441: outdata = 32'd50095;
			15442: outdata = 32'd50094;
			15443: outdata = 32'd50093;
			15444: outdata = 32'd50092;
			15445: outdata = 32'd50091;
			15446: outdata = 32'd50090;
			15447: outdata = 32'd50089;
			15448: outdata = 32'd50088;
			15449: outdata = 32'd50087;
			15450: outdata = 32'd50086;
			15451: outdata = 32'd50085;
			15452: outdata = 32'd50084;
			15453: outdata = 32'd50083;
			15454: outdata = 32'd50082;
			15455: outdata = 32'd50081;
			15456: outdata = 32'd50080;
			15457: outdata = 32'd50079;
			15458: outdata = 32'd50078;
			15459: outdata = 32'd50077;
			15460: outdata = 32'd50076;
			15461: outdata = 32'd50075;
			15462: outdata = 32'd50074;
			15463: outdata = 32'd50073;
			15464: outdata = 32'd50072;
			15465: outdata = 32'd50071;
			15466: outdata = 32'd50070;
			15467: outdata = 32'd50069;
			15468: outdata = 32'd50068;
			15469: outdata = 32'd50067;
			15470: outdata = 32'd50066;
			15471: outdata = 32'd50065;
			15472: outdata = 32'd50064;
			15473: outdata = 32'd50063;
			15474: outdata = 32'd50062;
			15475: outdata = 32'd50061;
			15476: outdata = 32'd50060;
			15477: outdata = 32'd50059;
			15478: outdata = 32'd50058;
			15479: outdata = 32'd50057;
			15480: outdata = 32'd50056;
			15481: outdata = 32'd50055;
			15482: outdata = 32'd50054;
			15483: outdata = 32'd50053;
			15484: outdata = 32'd50052;
			15485: outdata = 32'd50051;
			15486: outdata = 32'd50050;
			15487: outdata = 32'd50049;
			15488: outdata = 32'd50048;
			15489: outdata = 32'd50047;
			15490: outdata = 32'd50046;
			15491: outdata = 32'd50045;
			15492: outdata = 32'd50044;
			15493: outdata = 32'd50043;
			15494: outdata = 32'd50042;
			15495: outdata = 32'd50041;
			15496: outdata = 32'd50040;
			15497: outdata = 32'd50039;
			15498: outdata = 32'd50038;
			15499: outdata = 32'd50037;
			15500: outdata = 32'd50036;
			15501: outdata = 32'd50035;
			15502: outdata = 32'd50034;
			15503: outdata = 32'd50033;
			15504: outdata = 32'd50032;
			15505: outdata = 32'd50031;
			15506: outdata = 32'd50030;
			15507: outdata = 32'd50029;
			15508: outdata = 32'd50028;
			15509: outdata = 32'd50027;
			15510: outdata = 32'd50026;
			15511: outdata = 32'd50025;
			15512: outdata = 32'd50024;
			15513: outdata = 32'd50023;
			15514: outdata = 32'd50022;
			15515: outdata = 32'd50021;
			15516: outdata = 32'd50020;
			15517: outdata = 32'd50019;
			15518: outdata = 32'd50018;
			15519: outdata = 32'd50017;
			15520: outdata = 32'd50016;
			15521: outdata = 32'd50015;
			15522: outdata = 32'd50014;
			15523: outdata = 32'd50013;
			15524: outdata = 32'd50012;
			15525: outdata = 32'd50011;
			15526: outdata = 32'd50010;
			15527: outdata = 32'd50009;
			15528: outdata = 32'd50008;
			15529: outdata = 32'd50007;
			15530: outdata = 32'd50006;
			15531: outdata = 32'd50005;
			15532: outdata = 32'd50004;
			15533: outdata = 32'd50003;
			15534: outdata = 32'd50002;
			15535: outdata = 32'd50001;
			15536: outdata = 32'd50000;
			15537: outdata = 32'd49999;
			15538: outdata = 32'd49998;
			15539: outdata = 32'd49997;
			15540: outdata = 32'd49996;
			15541: outdata = 32'd49995;
			15542: outdata = 32'd49994;
			15543: outdata = 32'd49993;
			15544: outdata = 32'd49992;
			15545: outdata = 32'd49991;
			15546: outdata = 32'd49990;
			15547: outdata = 32'd49989;
			15548: outdata = 32'd49988;
			15549: outdata = 32'd49987;
			15550: outdata = 32'd49986;
			15551: outdata = 32'd49985;
			15552: outdata = 32'd49984;
			15553: outdata = 32'd49983;
			15554: outdata = 32'd49982;
			15555: outdata = 32'd49981;
			15556: outdata = 32'd49980;
			15557: outdata = 32'd49979;
			15558: outdata = 32'd49978;
			15559: outdata = 32'd49977;
			15560: outdata = 32'd49976;
			15561: outdata = 32'd49975;
			15562: outdata = 32'd49974;
			15563: outdata = 32'd49973;
			15564: outdata = 32'd49972;
			15565: outdata = 32'd49971;
			15566: outdata = 32'd49970;
			15567: outdata = 32'd49969;
			15568: outdata = 32'd49968;
			15569: outdata = 32'd49967;
			15570: outdata = 32'd49966;
			15571: outdata = 32'd49965;
			15572: outdata = 32'd49964;
			15573: outdata = 32'd49963;
			15574: outdata = 32'd49962;
			15575: outdata = 32'd49961;
			15576: outdata = 32'd49960;
			15577: outdata = 32'd49959;
			15578: outdata = 32'd49958;
			15579: outdata = 32'd49957;
			15580: outdata = 32'd49956;
			15581: outdata = 32'd49955;
			15582: outdata = 32'd49954;
			15583: outdata = 32'd49953;
			15584: outdata = 32'd49952;
			15585: outdata = 32'd49951;
			15586: outdata = 32'd49950;
			15587: outdata = 32'd49949;
			15588: outdata = 32'd49948;
			15589: outdata = 32'd49947;
			15590: outdata = 32'd49946;
			15591: outdata = 32'd49945;
			15592: outdata = 32'd49944;
			15593: outdata = 32'd49943;
			15594: outdata = 32'd49942;
			15595: outdata = 32'd49941;
			15596: outdata = 32'd49940;
			15597: outdata = 32'd49939;
			15598: outdata = 32'd49938;
			15599: outdata = 32'd49937;
			15600: outdata = 32'd49936;
			15601: outdata = 32'd49935;
			15602: outdata = 32'd49934;
			15603: outdata = 32'd49933;
			15604: outdata = 32'd49932;
			15605: outdata = 32'd49931;
			15606: outdata = 32'd49930;
			15607: outdata = 32'd49929;
			15608: outdata = 32'd49928;
			15609: outdata = 32'd49927;
			15610: outdata = 32'd49926;
			15611: outdata = 32'd49925;
			15612: outdata = 32'd49924;
			15613: outdata = 32'd49923;
			15614: outdata = 32'd49922;
			15615: outdata = 32'd49921;
			15616: outdata = 32'd49920;
			15617: outdata = 32'd49919;
			15618: outdata = 32'd49918;
			15619: outdata = 32'd49917;
			15620: outdata = 32'd49916;
			15621: outdata = 32'd49915;
			15622: outdata = 32'd49914;
			15623: outdata = 32'd49913;
			15624: outdata = 32'd49912;
			15625: outdata = 32'd49911;
			15626: outdata = 32'd49910;
			15627: outdata = 32'd49909;
			15628: outdata = 32'd49908;
			15629: outdata = 32'd49907;
			15630: outdata = 32'd49906;
			15631: outdata = 32'd49905;
			15632: outdata = 32'd49904;
			15633: outdata = 32'd49903;
			15634: outdata = 32'd49902;
			15635: outdata = 32'd49901;
			15636: outdata = 32'd49900;
			15637: outdata = 32'd49899;
			15638: outdata = 32'd49898;
			15639: outdata = 32'd49897;
			15640: outdata = 32'd49896;
			15641: outdata = 32'd49895;
			15642: outdata = 32'd49894;
			15643: outdata = 32'd49893;
			15644: outdata = 32'd49892;
			15645: outdata = 32'd49891;
			15646: outdata = 32'd49890;
			15647: outdata = 32'd49889;
			15648: outdata = 32'd49888;
			15649: outdata = 32'd49887;
			15650: outdata = 32'd49886;
			15651: outdata = 32'd49885;
			15652: outdata = 32'd49884;
			15653: outdata = 32'd49883;
			15654: outdata = 32'd49882;
			15655: outdata = 32'd49881;
			15656: outdata = 32'd49880;
			15657: outdata = 32'd49879;
			15658: outdata = 32'd49878;
			15659: outdata = 32'd49877;
			15660: outdata = 32'd49876;
			15661: outdata = 32'd49875;
			15662: outdata = 32'd49874;
			15663: outdata = 32'd49873;
			15664: outdata = 32'd49872;
			15665: outdata = 32'd49871;
			15666: outdata = 32'd49870;
			15667: outdata = 32'd49869;
			15668: outdata = 32'd49868;
			15669: outdata = 32'd49867;
			15670: outdata = 32'd49866;
			15671: outdata = 32'd49865;
			15672: outdata = 32'd49864;
			15673: outdata = 32'd49863;
			15674: outdata = 32'd49862;
			15675: outdata = 32'd49861;
			15676: outdata = 32'd49860;
			15677: outdata = 32'd49859;
			15678: outdata = 32'd49858;
			15679: outdata = 32'd49857;
			15680: outdata = 32'd49856;
			15681: outdata = 32'd49855;
			15682: outdata = 32'd49854;
			15683: outdata = 32'd49853;
			15684: outdata = 32'd49852;
			15685: outdata = 32'd49851;
			15686: outdata = 32'd49850;
			15687: outdata = 32'd49849;
			15688: outdata = 32'd49848;
			15689: outdata = 32'd49847;
			15690: outdata = 32'd49846;
			15691: outdata = 32'd49845;
			15692: outdata = 32'd49844;
			15693: outdata = 32'd49843;
			15694: outdata = 32'd49842;
			15695: outdata = 32'd49841;
			15696: outdata = 32'd49840;
			15697: outdata = 32'd49839;
			15698: outdata = 32'd49838;
			15699: outdata = 32'd49837;
			15700: outdata = 32'd49836;
			15701: outdata = 32'd49835;
			15702: outdata = 32'd49834;
			15703: outdata = 32'd49833;
			15704: outdata = 32'd49832;
			15705: outdata = 32'd49831;
			15706: outdata = 32'd49830;
			15707: outdata = 32'd49829;
			15708: outdata = 32'd49828;
			15709: outdata = 32'd49827;
			15710: outdata = 32'd49826;
			15711: outdata = 32'd49825;
			15712: outdata = 32'd49824;
			15713: outdata = 32'd49823;
			15714: outdata = 32'd49822;
			15715: outdata = 32'd49821;
			15716: outdata = 32'd49820;
			15717: outdata = 32'd49819;
			15718: outdata = 32'd49818;
			15719: outdata = 32'd49817;
			15720: outdata = 32'd49816;
			15721: outdata = 32'd49815;
			15722: outdata = 32'd49814;
			15723: outdata = 32'd49813;
			15724: outdata = 32'd49812;
			15725: outdata = 32'd49811;
			15726: outdata = 32'd49810;
			15727: outdata = 32'd49809;
			15728: outdata = 32'd49808;
			15729: outdata = 32'd49807;
			15730: outdata = 32'd49806;
			15731: outdata = 32'd49805;
			15732: outdata = 32'd49804;
			15733: outdata = 32'd49803;
			15734: outdata = 32'd49802;
			15735: outdata = 32'd49801;
			15736: outdata = 32'd49800;
			15737: outdata = 32'd49799;
			15738: outdata = 32'd49798;
			15739: outdata = 32'd49797;
			15740: outdata = 32'd49796;
			15741: outdata = 32'd49795;
			15742: outdata = 32'd49794;
			15743: outdata = 32'd49793;
			15744: outdata = 32'd49792;
			15745: outdata = 32'd49791;
			15746: outdata = 32'd49790;
			15747: outdata = 32'd49789;
			15748: outdata = 32'd49788;
			15749: outdata = 32'd49787;
			15750: outdata = 32'd49786;
			15751: outdata = 32'd49785;
			15752: outdata = 32'd49784;
			15753: outdata = 32'd49783;
			15754: outdata = 32'd49782;
			15755: outdata = 32'd49781;
			15756: outdata = 32'd49780;
			15757: outdata = 32'd49779;
			15758: outdata = 32'd49778;
			15759: outdata = 32'd49777;
			15760: outdata = 32'd49776;
			15761: outdata = 32'd49775;
			15762: outdata = 32'd49774;
			15763: outdata = 32'd49773;
			15764: outdata = 32'd49772;
			15765: outdata = 32'd49771;
			15766: outdata = 32'd49770;
			15767: outdata = 32'd49769;
			15768: outdata = 32'd49768;
			15769: outdata = 32'd49767;
			15770: outdata = 32'd49766;
			15771: outdata = 32'd49765;
			15772: outdata = 32'd49764;
			15773: outdata = 32'd49763;
			15774: outdata = 32'd49762;
			15775: outdata = 32'd49761;
			15776: outdata = 32'd49760;
			15777: outdata = 32'd49759;
			15778: outdata = 32'd49758;
			15779: outdata = 32'd49757;
			15780: outdata = 32'd49756;
			15781: outdata = 32'd49755;
			15782: outdata = 32'd49754;
			15783: outdata = 32'd49753;
			15784: outdata = 32'd49752;
			15785: outdata = 32'd49751;
			15786: outdata = 32'd49750;
			15787: outdata = 32'd49749;
			15788: outdata = 32'd49748;
			15789: outdata = 32'd49747;
			15790: outdata = 32'd49746;
			15791: outdata = 32'd49745;
			15792: outdata = 32'd49744;
			15793: outdata = 32'd49743;
			15794: outdata = 32'd49742;
			15795: outdata = 32'd49741;
			15796: outdata = 32'd49740;
			15797: outdata = 32'd49739;
			15798: outdata = 32'd49738;
			15799: outdata = 32'd49737;
			15800: outdata = 32'd49736;
			15801: outdata = 32'd49735;
			15802: outdata = 32'd49734;
			15803: outdata = 32'd49733;
			15804: outdata = 32'd49732;
			15805: outdata = 32'd49731;
			15806: outdata = 32'd49730;
			15807: outdata = 32'd49729;
			15808: outdata = 32'd49728;
			15809: outdata = 32'd49727;
			15810: outdata = 32'd49726;
			15811: outdata = 32'd49725;
			15812: outdata = 32'd49724;
			15813: outdata = 32'd49723;
			15814: outdata = 32'd49722;
			15815: outdata = 32'd49721;
			15816: outdata = 32'd49720;
			15817: outdata = 32'd49719;
			15818: outdata = 32'd49718;
			15819: outdata = 32'd49717;
			15820: outdata = 32'd49716;
			15821: outdata = 32'd49715;
			15822: outdata = 32'd49714;
			15823: outdata = 32'd49713;
			15824: outdata = 32'd49712;
			15825: outdata = 32'd49711;
			15826: outdata = 32'd49710;
			15827: outdata = 32'd49709;
			15828: outdata = 32'd49708;
			15829: outdata = 32'd49707;
			15830: outdata = 32'd49706;
			15831: outdata = 32'd49705;
			15832: outdata = 32'd49704;
			15833: outdata = 32'd49703;
			15834: outdata = 32'd49702;
			15835: outdata = 32'd49701;
			15836: outdata = 32'd49700;
			15837: outdata = 32'd49699;
			15838: outdata = 32'd49698;
			15839: outdata = 32'd49697;
			15840: outdata = 32'd49696;
			15841: outdata = 32'd49695;
			15842: outdata = 32'd49694;
			15843: outdata = 32'd49693;
			15844: outdata = 32'd49692;
			15845: outdata = 32'd49691;
			15846: outdata = 32'd49690;
			15847: outdata = 32'd49689;
			15848: outdata = 32'd49688;
			15849: outdata = 32'd49687;
			15850: outdata = 32'd49686;
			15851: outdata = 32'd49685;
			15852: outdata = 32'd49684;
			15853: outdata = 32'd49683;
			15854: outdata = 32'd49682;
			15855: outdata = 32'd49681;
			15856: outdata = 32'd49680;
			15857: outdata = 32'd49679;
			15858: outdata = 32'd49678;
			15859: outdata = 32'd49677;
			15860: outdata = 32'd49676;
			15861: outdata = 32'd49675;
			15862: outdata = 32'd49674;
			15863: outdata = 32'd49673;
			15864: outdata = 32'd49672;
			15865: outdata = 32'd49671;
			15866: outdata = 32'd49670;
			15867: outdata = 32'd49669;
			15868: outdata = 32'd49668;
			15869: outdata = 32'd49667;
			15870: outdata = 32'd49666;
			15871: outdata = 32'd49665;
			15872: outdata = 32'd49664;
			15873: outdata = 32'd49663;
			15874: outdata = 32'd49662;
			15875: outdata = 32'd49661;
			15876: outdata = 32'd49660;
			15877: outdata = 32'd49659;
			15878: outdata = 32'd49658;
			15879: outdata = 32'd49657;
			15880: outdata = 32'd49656;
			15881: outdata = 32'd49655;
			15882: outdata = 32'd49654;
			15883: outdata = 32'd49653;
			15884: outdata = 32'd49652;
			15885: outdata = 32'd49651;
			15886: outdata = 32'd49650;
			15887: outdata = 32'd49649;
			15888: outdata = 32'd49648;
			15889: outdata = 32'd49647;
			15890: outdata = 32'd49646;
			15891: outdata = 32'd49645;
			15892: outdata = 32'd49644;
			15893: outdata = 32'd49643;
			15894: outdata = 32'd49642;
			15895: outdata = 32'd49641;
			15896: outdata = 32'd49640;
			15897: outdata = 32'd49639;
			15898: outdata = 32'd49638;
			15899: outdata = 32'd49637;
			15900: outdata = 32'd49636;
			15901: outdata = 32'd49635;
			15902: outdata = 32'd49634;
			15903: outdata = 32'd49633;
			15904: outdata = 32'd49632;
			15905: outdata = 32'd49631;
			15906: outdata = 32'd49630;
			15907: outdata = 32'd49629;
			15908: outdata = 32'd49628;
			15909: outdata = 32'd49627;
			15910: outdata = 32'd49626;
			15911: outdata = 32'd49625;
			15912: outdata = 32'd49624;
			15913: outdata = 32'd49623;
			15914: outdata = 32'd49622;
			15915: outdata = 32'd49621;
			15916: outdata = 32'd49620;
			15917: outdata = 32'd49619;
			15918: outdata = 32'd49618;
			15919: outdata = 32'd49617;
			15920: outdata = 32'd49616;
			15921: outdata = 32'd49615;
			15922: outdata = 32'd49614;
			15923: outdata = 32'd49613;
			15924: outdata = 32'd49612;
			15925: outdata = 32'd49611;
			15926: outdata = 32'd49610;
			15927: outdata = 32'd49609;
			15928: outdata = 32'd49608;
			15929: outdata = 32'd49607;
			15930: outdata = 32'd49606;
			15931: outdata = 32'd49605;
			15932: outdata = 32'd49604;
			15933: outdata = 32'd49603;
			15934: outdata = 32'd49602;
			15935: outdata = 32'd49601;
			15936: outdata = 32'd49600;
			15937: outdata = 32'd49599;
			15938: outdata = 32'd49598;
			15939: outdata = 32'd49597;
			15940: outdata = 32'd49596;
			15941: outdata = 32'd49595;
			15942: outdata = 32'd49594;
			15943: outdata = 32'd49593;
			15944: outdata = 32'd49592;
			15945: outdata = 32'd49591;
			15946: outdata = 32'd49590;
			15947: outdata = 32'd49589;
			15948: outdata = 32'd49588;
			15949: outdata = 32'd49587;
			15950: outdata = 32'd49586;
			15951: outdata = 32'd49585;
			15952: outdata = 32'd49584;
			15953: outdata = 32'd49583;
			15954: outdata = 32'd49582;
			15955: outdata = 32'd49581;
			15956: outdata = 32'd49580;
			15957: outdata = 32'd49579;
			15958: outdata = 32'd49578;
			15959: outdata = 32'd49577;
			15960: outdata = 32'd49576;
			15961: outdata = 32'd49575;
			15962: outdata = 32'd49574;
			15963: outdata = 32'd49573;
			15964: outdata = 32'd49572;
			15965: outdata = 32'd49571;
			15966: outdata = 32'd49570;
			15967: outdata = 32'd49569;
			15968: outdata = 32'd49568;
			15969: outdata = 32'd49567;
			15970: outdata = 32'd49566;
			15971: outdata = 32'd49565;
			15972: outdata = 32'd49564;
			15973: outdata = 32'd49563;
			15974: outdata = 32'd49562;
			15975: outdata = 32'd49561;
			15976: outdata = 32'd49560;
			15977: outdata = 32'd49559;
			15978: outdata = 32'd49558;
			15979: outdata = 32'd49557;
			15980: outdata = 32'd49556;
			15981: outdata = 32'd49555;
			15982: outdata = 32'd49554;
			15983: outdata = 32'd49553;
			15984: outdata = 32'd49552;
			15985: outdata = 32'd49551;
			15986: outdata = 32'd49550;
			15987: outdata = 32'd49549;
			15988: outdata = 32'd49548;
			15989: outdata = 32'd49547;
			15990: outdata = 32'd49546;
			15991: outdata = 32'd49545;
			15992: outdata = 32'd49544;
			15993: outdata = 32'd49543;
			15994: outdata = 32'd49542;
			15995: outdata = 32'd49541;
			15996: outdata = 32'd49540;
			15997: outdata = 32'd49539;
			15998: outdata = 32'd49538;
			15999: outdata = 32'd49537;
			16000: outdata = 32'd49536;
			16001: outdata = 32'd49535;
			16002: outdata = 32'd49534;
			16003: outdata = 32'd49533;
			16004: outdata = 32'd49532;
			16005: outdata = 32'd49531;
			16006: outdata = 32'd49530;
			16007: outdata = 32'd49529;
			16008: outdata = 32'd49528;
			16009: outdata = 32'd49527;
			16010: outdata = 32'd49526;
			16011: outdata = 32'd49525;
			16012: outdata = 32'd49524;
			16013: outdata = 32'd49523;
			16014: outdata = 32'd49522;
			16015: outdata = 32'd49521;
			16016: outdata = 32'd49520;
			16017: outdata = 32'd49519;
			16018: outdata = 32'd49518;
			16019: outdata = 32'd49517;
			16020: outdata = 32'd49516;
			16021: outdata = 32'd49515;
			16022: outdata = 32'd49514;
			16023: outdata = 32'd49513;
			16024: outdata = 32'd49512;
			16025: outdata = 32'd49511;
			16026: outdata = 32'd49510;
			16027: outdata = 32'd49509;
			16028: outdata = 32'd49508;
			16029: outdata = 32'd49507;
			16030: outdata = 32'd49506;
			16031: outdata = 32'd49505;
			16032: outdata = 32'd49504;
			16033: outdata = 32'd49503;
			16034: outdata = 32'd49502;
			16035: outdata = 32'd49501;
			16036: outdata = 32'd49500;
			16037: outdata = 32'd49499;
			16038: outdata = 32'd49498;
			16039: outdata = 32'd49497;
			16040: outdata = 32'd49496;
			16041: outdata = 32'd49495;
			16042: outdata = 32'd49494;
			16043: outdata = 32'd49493;
			16044: outdata = 32'd49492;
			16045: outdata = 32'd49491;
			16046: outdata = 32'd49490;
			16047: outdata = 32'd49489;
			16048: outdata = 32'd49488;
			16049: outdata = 32'd49487;
			16050: outdata = 32'd49486;
			16051: outdata = 32'd49485;
			16052: outdata = 32'd49484;
			16053: outdata = 32'd49483;
			16054: outdata = 32'd49482;
			16055: outdata = 32'd49481;
			16056: outdata = 32'd49480;
			16057: outdata = 32'd49479;
			16058: outdata = 32'd49478;
			16059: outdata = 32'd49477;
			16060: outdata = 32'd49476;
			16061: outdata = 32'd49475;
			16062: outdata = 32'd49474;
			16063: outdata = 32'd49473;
			16064: outdata = 32'd49472;
			16065: outdata = 32'd49471;
			16066: outdata = 32'd49470;
			16067: outdata = 32'd49469;
			16068: outdata = 32'd49468;
			16069: outdata = 32'd49467;
			16070: outdata = 32'd49466;
			16071: outdata = 32'd49465;
			16072: outdata = 32'd49464;
			16073: outdata = 32'd49463;
			16074: outdata = 32'd49462;
			16075: outdata = 32'd49461;
			16076: outdata = 32'd49460;
			16077: outdata = 32'd49459;
			16078: outdata = 32'd49458;
			16079: outdata = 32'd49457;
			16080: outdata = 32'd49456;
			16081: outdata = 32'd49455;
			16082: outdata = 32'd49454;
			16083: outdata = 32'd49453;
			16084: outdata = 32'd49452;
			16085: outdata = 32'd49451;
			16086: outdata = 32'd49450;
			16087: outdata = 32'd49449;
			16088: outdata = 32'd49448;
			16089: outdata = 32'd49447;
			16090: outdata = 32'd49446;
			16091: outdata = 32'd49445;
			16092: outdata = 32'd49444;
			16093: outdata = 32'd49443;
			16094: outdata = 32'd49442;
			16095: outdata = 32'd49441;
			16096: outdata = 32'd49440;
			16097: outdata = 32'd49439;
			16098: outdata = 32'd49438;
			16099: outdata = 32'd49437;
			16100: outdata = 32'd49436;
			16101: outdata = 32'd49435;
			16102: outdata = 32'd49434;
			16103: outdata = 32'd49433;
			16104: outdata = 32'd49432;
			16105: outdata = 32'd49431;
			16106: outdata = 32'd49430;
			16107: outdata = 32'd49429;
			16108: outdata = 32'd49428;
			16109: outdata = 32'd49427;
			16110: outdata = 32'd49426;
			16111: outdata = 32'd49425;
			16112: outdata = 32'd49424;
			16113: outdata = 32'd49423;
			16114: outdata = 32'd49422;
			16115: outdata = 32'd49421;
			16116: outdata = 32'd49420;
			16117: outdata = 32'd49419;
			16118: outdata = 32'd49418;
			16119: outdata = 32'd49417;
			16120: outdata = 32'd49416;
			16121: outdata = 32'd49415;
			16122: outdata = 32'd49414;
			16123: outdata = 32'd49413;
			16124: outdata = 32'd49412;
			16125: outdata = 32'd49411;
			16126: outdata = 32'd49410;
			16127: outdata = 32'd49409;
			16128: outdata = 32'd49408;
			16129: outdata = 32'd49407;
			16130: outdata = 32'd49406;
			16131: outdata = 32'd49405;
			16132: outdata = 32'd49404;
			16133: outdata = 32'd49403;
			16134: outdata = 32'd49402;
			16135: outdata = 32'd49401;
			16136: outdata = 32'd49400;
			16137: outdata = 32'd49399;
			16138: outdata = 32'd49398;
			16139: outdata = 32'd49397;
			16140: outdata = 32'd49396;
			16141: outdata = 32'd49395;
			16142: outdata = 32'd49394;
			16143: outdata = 32'd49393;
			16144: outdata = 32'd49392;
			16145: outdata = 32'd49391;
			16146: outdata = 32'd49390;
			16147: outdata = 32'd49389;
			16148: outdata = 32'd49388;
			16149: outdata = 32'd49387;
			16150: outdata = 32'd49386;
			16151: outdata = 32'd49385;
			16152: outdata = 32'd49384;
			16153: outdata = 32'd49383;
			16154: outdata = 32'd49382;
			16155: outdata = 32'd49381;
			16156: outdata = 32'd49380;
			16157: outdata = 32'd49379;
			16158: outdata = 32'd49378;
			16159: outdata = 32'd49377;
			16160: outdata = 32'd49376;
			16161: outdata = 32'd49375;
			16162: outdata = 32'd49374;
			16163: outdata = 32'd49373;
			16164: outdata = 32'd49372;
			16165: outdata = 32'd49371;
			16166: outdata = 32'd49370;
			16167: outdata = 32'd49369;
			16168: outdata = 32'd49368;
			16169: outdata = 32'd49367;
			16170: outdata = 32'd49366;
			16171: outdata = 32'd49365;
			16172: outdata = 32'd49364;
			16173: outdata = 32'd49363;
			16174: outdata = 32'd49362;
			16175: outdata = 32'd49361;
			16176: outdata = 32'd49360;
			16177: outdata = 32'd49359;
			16178: outdata = 32'd49358;
			16179: outdata = 32'd49357;
			16180: outdata = 32'd49356;
			16181: outdata = 32'd49355;
			16182: outdata = 32'd49354;
			16183: outdata = 32'd49353;
			16184: outdata = 32'd49352;
			16185: outdata = 32'd49351;
			16186: outdata = 32'd49350;
			16187: outdata = 32'd49349;
			16188: outdata = 32'd49348;
			16189: outdata = 32'd49347;
			16190: outdata = 32'd49346;
			16191: outdata = 32'd49345;
			16192: outdata = 32'd49344;
			16193: outdata = 32'd49343;
			16194: outdata = 32'd49342;
			16195: outdata = 32'd49341;
			16196: outdata = 32'd49340;
			16197: outdata = 32'd49339;
			16198: outdata = 32'd49338;
			16199: outdata = 32'd49337;
			16200: outdata = 32'd49336;
			16201: outdata = 32'd49335;
			16202: outdata = 32'd49334;
			16203: outdata = 32'd49333;
			16204: outdata = 32'd49332;
			16205: outdata = 32'd49331;
			16206: outdata = 32'd49330;
			16207: outdata = 32'd49329;
			16208: outdata = 32'd49328;
			16209: outdata = 32'd49327;
			16210: outdata = 32'd49326;
			16211: outdata = 32'd49325;
			16212: outdata = 32'd49324;
			16213: outdata = 32'd49323;
			16214: outdata = 32'd49322;
			16215: outdata = 32'd49321;
			16216: outdata = 32'd49320;
			16217: outdata = 32'd49319;
			16218: outdata = 32'd49318;
			16219: outdata = 32'd49317;
			16220: outdata = 32'd49316;
			16221: outdata = 32'd49315;
			16222: outdata = 32'd49314;
			16223: outdata = 32'd49313;
			16224: outdata = 32'd49312;
			16225: outdata = 32'd49311;
			16226: outdata = 32'd49310;
			16227: outdata = 32'd49309;
			16228: outdata = 32'd49308;
			16229: outdata = 32'd49307;
			16230: outdata = 32'd49306;
			16231: outdata = 32'd49305;
			16232: outdata = 32'd49304;
			16233: outdata = 32'd49303;
			16234: outdata = 32'd49302;
			16235: outdata = 32'd49301;
			16236: outdata = 32'd49300;
			16237: outdata = 32'd49299;
			16238: outdata = 32'd49298;
			16239: outdata = 32'd49297;
			16240: outdata = 32'd49296;
			16241: outdata = 32'd49295;
			16242: outdata = 32'd49294;
			16243: outdata = 32'd49293;
			16244: outdata = 32'd49292;
			16245: outdata = 32'd49291;
			16246: outdata = 32'd49290;
			16247: outdata = 32'd49289;
			16248: outdata = 32'd49288;
			16249: outdata = 32'd49287;
			16250: outdata = 32'd49286;
			16251: outdata = 32'd49285;
			16252: outdata = 32'd49284;
			16253: outdata = 32'd49283;
			16254: outdata = 32'd49282;
			16255: outdata = 32'd49281;
			16256: outdata = 32'd49280;
			16257: outdata = 32'd49279;
			16258: outdata = 32'd49278;
			16259: outdata = 32'd49277;
			16260: outdata = 32'd49276;
			16261: outdata = 32'd49275;
			16262: outdata = 32'd49274;
			16263: outdata = 32'd49273;
			16264: outdata = 32'd49272;
			16265: outdata = 32'd49271;
			16266: outdata = 32'd49270;
			16267: outdata = 32'd49269;
			16268: outdata = 32'd49268;
			16269: outdata = 32'd49267;
			16270: outdata = 32'd49266;
			16271: outdata = 32'd49265;
			16272: outdata = 32'd49264;
			16273: outdata = 32'd49263;
			16274: outdata = 32'd49262;
			16275: outdata = 32'd49261;
			16276: outdata = 32'd49260;
			16277: outdata = 32'd49259;
			16278: outdata = 32'd49258;
			16279: outdata = 32'd49257;
			16280: outdata = 32'd49256;
			16281: outdata = 32'd49255;
			16282: outdata = 32'd49254;
			16283: outdata = 32'd49253;
			16284: outdata = 32'd49252;
			16285: outdata = 32'd49251;
			16286: outdata = 32'd49250;
			16287: outdata = 32'd49249;
			16288: outdata = 32'd49248;
			16289: outdata = 32'd49247;
			16290: outdata = 32'd49246;
			16291: outdata = 32'd49245;
			16292: outdata = 32'd49244;
			16293: outdata = 32'd49243;
			16294: outdata = 32'd49242;
			16295: outdata = 32'd49241;
			16296: outdata = 32'd49240;
			16297: outdata = 32'd49239;
			16298: outdata = 32'd49238;
			16299: outdata = 32'd49237;
			16300: outdata = 32'd49236;
			16301: outdata = 32'd49235;
			16302: outdata = 32'd49234;
			16303: outdata = 32'd49233;
			16304: outdata = 32'd49232;
			16305: outdata = 32'd49231;
			16306: outdata = 32'd49230;
			16307: outdata = 32'd49229;
			16308: outdata = 32'd49228;
			16309: outdata = 32'd49227;
			16310: outdata = 32'd49226;
			16311: outdata = 32'd49225;
			16312: outdata = 32'd49224;
			16313: outdata = 32'd49223;
			16314: outdata = 32'd49222;
			16315: outdata = 32'd49221;
			16316: outdata = 32'd49220;
			16317: outdata = 32'd49219;
			16318: outdata = 32'd49218;
			16319: outdata = 32'd49217;
			16320: outdata = 32'd49216;
			16321: outdata = 32'd49215;
			16322: outdata = 32'd49214;
			16323: outdata = 32'd49213;
			16324: outdata = 32'd49212;
			16325: outdata = 32'd49211;
			16326: outdata = 32'd49210;
			16327: outdata = 32'd49209;
			16328: outdata = 32'd49208;
			16329: outdata = 32'd49207;
			16330: outdata = 32'd49206;
			16331: outdata = 32'd49205;
			16332: outdata = 32'd49204;
			16333: outdata = 32'd49203;
			16334: outdata = 32'd49202;
			16335: outdata = 32'd49201;
			16336: outdata = 32'd49200;
			16337: outdata = 32'd49199;
			16338: outdata = 32'd49198;
			16339: outdata = 32'd49197;
			16340: outdata = 32'd49196;
			16341: outdata = 32'd49195;
			16342: outdata = 32'd49194;
			16343: outdata = 32'd49193;
			16344: outdata = 32'd49192;
			16345: outdata = 32'd49191;
			16346: outdata = 32'd49190;
			16347: outdata = 32'd49189;
			16348: outdata = 32'd49188;
			16349: outdata = 32'd49187;
			16350: outdata = 32'd49186;
			16351: outdata = 32'd49185;
			16352: outdata = 32'd49184;
			16353: outdata = 32'd49183;
			16354: outdata = 32'd49182;
			16355: outdata = 32'd49181;
			16356: outdata = 32'd49180;
			16357: outdata = 32'd49179;
			16358: outdata = 32'd49178;
			16359: outdata = 32'd49177;
			16360: outdata = 32'd49176;
			16361: outdata = 32'd49175;
			16362: outdata = 32'd49174;
			16363: outdata = 32'd49173;
			16364: outdata = 32'd49172;
			16365: outdata = 32'd49171;
			16366: outdata = 32'd49170;
			16367: outdata = 32'd49169;
			16368: outdata = 32'd49168;
			16369: outdata = 32'd49167;
			16370: outdata = 32'd49166;
			16371: outdata = 32'd49165;
			16372: outdata = 32'd49164;
			16373: outdata = 32'd49163;
			16374: outdata = 32'd49162;
			16375: outdata = 32'd49161;
			16376: outdata = 32'd49160;
			16377: outdata = 32'd49159;
			16378: outdata = 32'd49158;
			16379: outdata = 32'd49157;
			16380: outdata = 32'd49156;
			16381: outdata = 32'd49155;
			16382: outdata = 32'd49154;
			16383: outdata = 32'd49153;
			16384: outdata = 32'd49152;
			16385: outdata = 32'd49151;
			16386: outdata = 32'd49150;
			16387: outdata = 32'd49149;
			16388: outdata = 32'd49148;
			16389: outdata = 32'd49147;
			16390: outdata = 32'd49146;
			16391: outdata = 32'd49145;
			16392: outdata = 32'd49144;
			16393: outdata = 32'd49143;
			16394: outdata = 32'd49142;
			16395: outdata = 32'd49141;
			16396: outdata = 32'd49140;
			16397: outdata = 32'd49139;
			16398: outdata = 32'd49138;
			16399: outdata = 32'd49137;
			16400: outdata = 32'd49136;
			16401: outdata = 32'd49135;
			16402: outdata = 32'd49134;
			16403: outdata = 32'd49133;
			16404: outdata = 32'd49132;
			16405: outdata = 32'd49131;
			16406: outdata = 32'd49130;
			16407: outdata = 32'd49129;
			16408: outdata = 32'd49128;
			16409: outdata = 32'd49127;
			16410: outdata = 32'd49126;
			16411: outdata = 32'd49125;
			16412: outdata = 32'd49124;
			16413: outdata = 32'd49123;
			16414: outdata = 32'd49122;
			16415: outdata = 32'd49121;
			16416: outdata = 32'd49120;
			16417: outdata = 32'd49119;
			16418: outdata = 32'd49118;
			16419: outdata = 32'd49117;
			16420: outdata = 32'd49116;
			16421: outdata = 32'd49115;
			16422: outdata = 32'd49114;
			16423: outdata = 32'd49113;
			16424: outdata = 32'd49112;
			16425: outdata = 32'd49111;
			16426: outdata = 32'd49110;
			16427: outdata = 32'd49109;
			16428: outdata = 32'd49108;
			16429: outdata = 32'd49107;
			16430: outdata = 32'd49106;
			16431: outdata = 32'd49105;
			16432: outdata = 32'd49104;
			16433: outdata = 32'd49103;
			16434: outdata = 32'd49102;
			16435: outdata = 32'd49101;
			16436: outdata = 32'd49100;
			16437: outdata = 32'd49099;
			16438: outdata = 32'd49098;
			16439: outdata = 32'd49097;
			16440: outdata = 32'd49096;
			16441: outdata = 32'd49095;
			16442: outdata = 32'd49094;
			16443: outdata = 32'd49093;
			16444: outdata = 32'd49092;
			16445: outdata = 32'd49091;
			16446: outdata = 32'd49090;
			16447: outdata = 32'd49089;
			16448: outdata = 32'd49088;
			16449: outdata = 32'd49087;
			16450: outdata = 32'd49086;
			16451: outdata = 32'd49085;
			16452: outdata = 32'd49084;
			16453: outdata = 32'd49083;
			16454: outdata = 32'd49082;
			16455: outdata = 32'd49081;
			16456: outdata = 32'd49080;
			16457: outdata = 32'd49079;
			16458: outdata = 32'd49078;
			16459: outdata = 32'd49077;
			16460: outdata = 32'd49076;
			16461: outdata = 32'd49075;
			16462: outdata = 32'd49074;
			16463: outdata = 32'd49073;
			16464: outdata = 32'd49072;
			16465: outdata = 32'd49071;
			16466: outdata = 32'd49070;
			16467: outdata = 32'd49069;
			16468: outdata = 32'd49068;
			16469: outdata = 32'd49067;
			16470: outdata = 32'd49066;
			16471: outdata = 32'd49065;
			16472: outdata = 32'd49064;
			16473: outdata = 32'd49063;
			16474: outdata = 32'd49062;
			16475: outdata = 32'd49061;
			16476: outdata = 32'd49060;
			16477: outdata = 32'd49059;
			16478: outdata = 32'd49058;
			16479: outdata = 32'd49057;
			16480: outdata = 32'd49056;
			16481: outdata = 32'd49055;
			16482: outdata = 32'd49054;
			16483: outdata = 32'd49053;
			16484: outdata = 32'd49052;
			16485: outdata = 32'd49051;
			16486: outdata = 32'd49050;
			16487: outdata = 32'd49049;
			16488: outdata = 32'd49048;
			16489: outdata = 32'd49047;
			16490: outdata = 32'd49046;
			16491: outdata = 32'd49045;
			16492: outdata = 32'd49044;
			16493: outdata = 32'd49043;
			16494: outdata = 32'd49042;
			16495: outdata = 32'd49041;
			16496: outdata = 32'd49040;
			16497: outdata = 32'd49039;
			16498: outdata = 32'd49038;
			16499: outdata = 32'd49037;
			16500: outdata = 32'd49036;
			16501: outdata = 32'd49035;
			16502: outdata = 32'd49034;
			16503: outdata = 32'd49033;
			16504: outdata = 32'd49032;
			16505: outdata = 32'd49031;
			16506: outdata = 32'd49030;
			16507: outdata = 32'd49029;
			16508: outdata = 32'd49028;
			16509: outdata = 32'd49027;
			16510: outdata = 32'd49026;
			16511: outdata = 32'd49025;
			16512: outdata = 32'd49024;
			16513: outdata = 32'd49023;
			16514: outdata = 32'd49022;
			16515: outdata = 32'd49021;
			16516: outdata = 32'd49020;
			16517: outdata = 32'd49019;
			16518: outdata = 32'd49018;
			16519: outdata = 32'd49017;
			16520: outdata = 32'd49016;
			16521: outdata = 32'd49015;
			16522: outdata = 32'd49014;
			16523: outdata = 32'd49013;
			16524: outdata = 32'd49012;
			16525: outdata = 32'd49011;
			16526: outdata = 32'd49010;
			16527: outdata = 32'd49009;
			16528: outdata = 32'd49008;
			16529: outdata = 32'd49007;
			16530: outdata = 32'd49006;
			16531: outdata = 32'd49005;
			16532: outdata = 32'd49004;
			16533: outdata = 32'd49003;
			16534: outdata = 32'd49002;
			16535: outdata = 32'd49001;
			16536: outdata = 32'd49000;
			16537: outdata = 32'd48999;
			16538: outdata = 32'd48998;
			16539: outdata = 32'd48997;
			16540: outdata = 32'd48996;
			16541: outdata = 32'd48995;
			16542: outdata = 32'd48994;
			16543: outdata = 32'd48993;
			16544: outdata = 32'd48992;
			16545: outdata = 32'd48991;
			16546: outdata = 32'd48990;
			16547: outdata = 32'd48989;
			16548: outdata = 32'd48988;
			16549: outdata = 32'd48987;
			16550: outdata = 32'd48986;
			16551: outdata = 32'd48985;
			16552: outdata = 32'd48984;
			16553: outdata = 32'd48983;
			16554: outdata = 32'd48982;
			16555: outdata = 32'd48981;
			16556: outdata = 32'd48980;
			16557: outdata = 32'd48979;
			16558: outdata = 32'd48978;
			16559: outdata = 32'd48977;
			16560: outdata = 32'd48976;
			16561: outdata = 32'd48975;
			16562: outdata = 32'd48974;
			16563: outdata = 32'd48973;
			16564: outdata = 32'd48972;
			16565: outdata = 32'd48971;
			16566: outdata = 32'd48970;
			16567: outdata = 32'd48969;
			16568: outdata = 32'd48968;
			16569: outdata = 32'd48967;
			16570: outdata = 32'd48966;
			16571: outdata = 32'd48965;
			16572: outdata = 32'd48964;
			16573: outdata = 32'd48963;
			16574: outdata = 32'd48962;
			16575: outdata = 32'd48961;
			16576: outdata = 32'd48960;
			16577: outdata = 32'd48959;
			16578: outdata = 32'd48958;
			16579: outdata = 32'd48957;
			16580: outdata = 32'd48956;
			16581: outdata = 32'd48955;
			16582: outdata = 32'd48954;
			16583: outdata = 32'd48953;
			16584: outdata = 32'd48952;
			16585: outdata = 32'd48951;
			16586: outdata = 32'd48950;
			16587: outdata = 32'd48949;
			16588: outdata = 32'd48948;
			16589: outdata = 32'd48947;
			16590: outdata = 32'd48946;
			16591: outdata = 32'd48945;
			16592: outdata = 32'd48944;
			16593: outdata = 32'd48943;
			16594: outdata = 32'd48942;
			16595: outdata = 32'd48941;
			16596: outdata = 32'd48940;
			16597: outdata = 32'd48939;
			16598: outdata = 32'd48938;
			16599: outdata = 32'd48937;
			16600: outdata = 32'd48936;
			16601: outdata = 32'd48935;
			16602: outdata = 32'd48934;
			16603: outdata = 32'd48933;
			16604: outdata = 32'd48932;
			16605: outdata = 32'd48931;
			16606: outdata = 32'd48930;
			16607: outdata = 32'd48929;
			16608: outdata = 32'd48928;
			16609: outdata = 32'd48927;
			16610: outdata = 32'd48926;
			16611: outdata = 32'd48925;
			16612: outdata = 32'd48924;
			16613: outdata = 32'd48923;
			16614: outdata = 32'd48922;
			16615: outdata = 32'd48921;
			16616: outdata = 32'd48920;
			16617: outdata = 32'd48919;
			16618: outdata = 32'd48918;
			16619: outdata = 32'd48917;
			16620: outdata = 32'd48916;
			16621: outdata = 32'd48915;
			16622: outdata = 32'd48914;
			16623: outdata = 32'd48913;
			16624: outdata = 32'd48912;
			16625: outdata = 32'd48911;
			16626: outdata = 32'd48910;
			16627: outdata = 32'd48909;
			16628: outdata = 32'd48908;
			16629: outdata = 32'd48907;
			16630: outdata = 32'd48906;
			16631: outdata = 32'd48905;
			16632: outdata = 32'd48904;
			16633: outdata = 32'd48903;
			16634: outdata = 32'd48902;
			16635: outdata = 32'd48901;
			16636: outdata = 32'd48900;
			16637: outdata = 32'd48899;
			16638: outdata = 32'd48898;
			16639: outdata = 32'd48897;
			16640: outdata = 32'd48896;
			16641: outdata = 32'd48895;
			16642: outdata = 32'd48894;
			16643: outdata = 32'd48893;
			16644: outdata = 32'd48892;
			16645: outdata = 32'd48891;
			16646: outdata = 32'd48890;
			16647: outdata = 32'd48889;
			16648: outdata = 32'd48888;
			16649: outdata = 32'd48887;
			16650: outdata = 32'd48886;
			16651: outdata = 32'd48885;
			16652: outdata = 32'd48884;
			16653: outdata = 32'd48883;
			16654: outdata = 32'd48882;
			16655: outdata = 32'd48881;
			16656: outdata = 32'd48880;
			16657: outdata = 32'd48879;
			16658: outdata = 32'd48878;
			16659: outdata = 32'd48877;
			16660: outdata = 32'd48876;
			16661: outdata = 32'd48875;
			16662: outdata = 32'd48874;
			16663: outdata = 32'd48873;
			16664: outdata = 32'd48872;
			16665: outdata = 32'd48871;
			16666: outdata = 32'd48870;
			16667: outdata = 32'd48869;
			16668: outdata = 32'd48868;
			16669: outdata = 32'd48867;
			16670: outdata = 32'd48866;
			16671: outdata = 32'd48865;
			16672: outdata = 32'd48864;
			16673: outdata = 32'd48863;
			16674: outdata = 32'd48862;
			16675: outdata = 32'd48861;
			16676: outdata = 32'd48860;
			16677: outdata = 32'd48859;
			16678: outdata = 32'd48858;
			16679: outdata = 32'd48857;
			16680: outdata = 32'd48856;
			16681: outdata = 32'd48855;
			16682: outdata = 32'd48854;
			16683: outdata = 32'd48853;
			16684: outdata = 32'd48852;
			16685: outdata = 32'd48851;
			16686: outdata = 32'd48850;
			16687: outdata = 32'd48849;
			16688: outdata = 32'd48848;
			16689: outdata = 32'd48847;
			16690: outdata = 32'd48846;
			16691: outdata = 32'd48845;
			16692: outdata = 32'd48844;
			16693: outdata = 32'd48843;
			16694: outdata = 32'd48842;
			16695: outdata = 32'd48841;
			16696: outdata = 32'd48840;
			16697: outdata = 32'd48839;
			16698: outdata = 32'd48838;
			16699: outdata = 32'd48837;
			16700: outdata = 32'd48836;
			16701: outdata = 32'd48835;
			16702: outdata = 32'd48834;
			16703: outdata = 32'd48833;
			16704: outdata = 32'd48832;
			16705: outdata = 32'd48831;
			16706: outdata = 32'd48830;
			16707: outdata = 32'd48829;
			16708: outdata = 32'd48828;
			16709: outdata = 32'd48827;
			16710: outdata = 32'd48826;
			16711: outdata = 32'd48825;
			16712: outdata = 32'd48824;
			16713: outdata = 32'd48823;
			16714: outdata = 32'd48822;
			16715: outdata = 32'd48821;
			16716: outdata = 32'd48820;
			16717: outdata = 32'd48819;
			16718: outdata = 32'd48818;
			16719: outdata = 32'd48817;
			16720: outdata = 32'd48816;
			16721: outdata = 32'd48815;
			16722: outdata = 32'd48814;
			16723: outdata = 32'd48813;
			16724: outdata = 32'd48812;
			16725: outdata = 32'd48811;
			16726: outdata = 32'd48810;
			16727: outdata = 32'd48809;
			16728: outdata = 32'd48808;
			16729: outdata = 32'd48807;
			16730: outdata = 32'd48806;
			16731: outdata = 32'd48805;
			16732: outdata = 32'd48804;
			16733: outdata = 32'd48803;
			16734: outdata = 32'd48802;
			16735: outdata = 32'd48801;
			16736: outdata = 32'd48800;
			16737: outdata = 32'd48799;
			16738: outdata = 32'd48798;
			16739: outdata = 32'd48797;
			16740: outdata = 32'd48796;
			16741: outdata = 32'd48795;
			16742: outdata = 32'd48794;
			16743: outdata = 32'd48793;
			16744: outdata = 32'd48792;
			16745: outdata = 32'd48791;
			16746: outdata = 32'd48790;
			16747: outdata = 32'd48789;
			16748: outdata = 32'd48788;
			16749: outdata = 32'd48787;
			16750: outdata = 32'd48786;
			16751: outdata = 32'd48785;
			16752: outdata = 32'd48784;
			16753: outdata = 32'd48783;
			16754: outdata = 32'd48782;
			16755: outdata = 32'd48781;
			16756: outdata = 32'd48780;
			16757: outdata = 32'd48779;
			16758: outdata = 32'd48778;
			16759: outdata = 32'd48777;
			16760: outdata = 32'd48776;
			16761: outdata = 32'd48775;
			16762: outdata = 32'd48774;
			16763: outdata = 32'd48773;
			16764: outdata = 32'd48772;
			16765: outdata = 32'd48771;
			16766: outdata = 32'd48770;
			16767: outdata = 32'd48769;
			16768: outdata = 32'd48768;
			16769: outdata = 32'd48767;
			16770: outdata = 32'd48766;
			16771: outdata = 32'd48765;
			16772: outdata = 32'd48764;
			16773: outdata = 32'd48763;
			16774: outdata = 32'd48762;
			16775: outdata = 32'd48761;
			16776: outdata = 32'd48760;
			16777: outdata = 32'd48759;
			16778: outdata = 32'd48758;
			16779: outdata = 32'd48757;
			16780: outdata = 32'd48756;
			16781: outdata = 32'd48755;
			16782: outdata = 32'd48754;
			16783: outdata = 32'd48753;
			16784: outdata = 32'd48752;
			16785: outdata = 32'd48751;
			16786: outdata = 32'd48750;
			16787: outdata = 32'd48749;
			16788: outdata = 32'd48748;
			16789: outdata = 32'd48747;
			16790: outdata = 32'd48746;
			16791: outdata = 32'd48745;
			16792: outdata = 32'd48744;
			16793: outdata = 32'd48743;
			16794: outdata = 32'd48742;
			16795: outdata = 32'd48741;
			16796: outdata = 32'd48740;
			16797: outdata = 32'd48739;
			16798: outdata = 32'd48738;
			16799: outdata = 32'd48737;
			16800: outdata = 32'd48736;
			16801: outdata = 32'd48735;
			16802: outdata = 32'd48734;
			16803: outdata = 32'd48733;
			16804: outdata = 32'd48732;
			16805: outdata = 32'd48731;
			16806: outdata = 32'd48730;
			16807: outdata = 32'd48729;
			16808: outdata = 32'd48728;
			16809: outdata = 32'd48727;
			16810: outdata = 32'd48726;
			16811: outdata = 32'd48725;
			16812: outdata = 32'd48724;
			16813: outdata = 32'd48723;
			16814: outdata = 32'd48722;
			16815: outdata = 32'd48721;
			16816: outdata = 32'd48720;
			16817: outdata = 32'd48719;
			16818: outdata = 32'd48718;
			16819: outdata = 32'd48717;
			16820: outdata = 32'd48716;
			16821: outdata = 32'd48715;
			16822: outdata = 32'd48714;
			16823: outdata = 32'd48713;
			16824: outdata = 32'd48712;
			16825: outdata = 32'd48711;
			16826: outdata = 32'd48710;
			16827: outdata = 32'd48709;
			16828: outdata = 32'd48708;
			16829: outdata = 32'd48707;
			16830: outdata = 32'd48706;
			16831: outdata = 32'd48705;
			16832: outdata = 32'd48704;
			16833: outdata = 32'd48703;
			16834: outdata = 32'd48702;
			16835: outdata = 32'd48701;
			16836: outdata = 32'd48700;
			16837: outdata = 32'd48699;
			16838: outdata = 32'd48698;
			16839: outdata = 32'd48697;
			16840: outdata = 32'd48696;
			16841: outdata = 32'd48695;
			16842: outdata = 32'd48694;
			16843: outdata = 32'd48693;
			16844: outdata = 32'd48692;
			16845: outdata = 32'd48691;
			16846: outdata = 32'd48690;
			16847: outdata = 32'd48689;
			16848: outdata = 32'd48688;
			16849: outdata = 32'd48687;
			16850: outdata = 32'd48686;
			16851: outdata = 32'd48685;
			16852: outdata = 32'd48684;
			16853: outdata = 32'd48683;
			16854: outdata = 32'd48682;
			16855: outdata = 32'd48681;
			16856: outdata = 32'd48680;
			16857: outdata = 32'd48679;
			16858: outdata = 32'd48678;
			16859: outdata = 32'd48677;
			16860: outdata = 32'd48676;
			16861: outdata = 32'd48675;
			16862: outdata = 32'd48674;
			16863: outdata = 32'd48673;
			16864: outdata = 32'd48672;
			16865: outdata = 32'd48671;
			16866: outdata = 32'd48670;
			16867: outdata = 32'd48669;
			16868: outdata = 32'd48668;
			16869: outdata = 32'd48667;
			16870: outdata = 32'd48666;
			16871: outdata = 32'd48665;
			16872: outdata = 32'd48664;
			16873: outdata = 32'd48663;
			16874: outdata = 32'd48662;
			16875: outdata = 32'd48661;
			16876: outdata = 32'd48660;
			16877: outdata = 32'd48659;
			16878: outdata = 32'd48658;
			16879: outdata = 32'd48657;
			16880: outdata = 32'd48656;
			16881: outdata = 32'd48655;
			16882: outdata = 32'd48654;
			16883: outdata = 32'd48653;
			16884: outdata = 32'd48652;
			16885: outdata = 32'd48651;
			16886: outdata = 32'd48650;
			16887: outdata = 32'd48649;
			16888: outdata = 32'd48648;
			16889: outdata = 32'd48647;
			16890: outdata = 32'd48646;
			16891: outdata = 32'd48645;
			16892: outdata = 32'd48644;
			16893: outdata = 32'd48643;
			16894: outdata = 32'd48642;
			16895: outdata = 32'd48641;
			16896: outdata = 32'd48640;
			16897: outdata = 32'd48639;
			16898: outdata = 32'd48638;
			16899: outdata = 32'd48637;
			16900: outdata = 32'd48636;
			16901: outdata = 32'd48635;
			16902: outdata = 32'd48634;
			16903: outdata = 32'd48633;
			16904: outdata = 32'd48632;
			16905: outdata = 32'd48631;
			16906: outdata = 32'd48630;
			16907: outdata = 32'd48629;
			16908: outdata = 32'd48628;
			16909: outdata = 32'd48627;
			16910: outdata = 32'd48626;
			16911: outdata = 32'd48625;
			16912: outdata = 32'd48624;
			16913: outdata = 32'd48623;
			16914: outdata = 32'd48622;
			16915: outdata = 32'd48621;
			16916: outdata = 32'd48620;
			16917: outdata = 32'd48619;
			16918: outdata = 32'd48618;
			16919: outdata = 32'd48617;
			16920: outdata = 32'd48616;
			16921: outdata = 32'd48615;
			16922: outdata = 32'd48614;
			16923: outdata = 32'd48613;
			16924: outdata = 32'd48612;
			16925: outdata = 32'd48611;
			16926: outdata = 32'd48610;
			16927: outdata = 32'd48609;
			16928: outdata = 32'd48608;
			16929: outdata = 32'd48607;
			16930: outdata = 32'd48606;
			16931: outdata = 32'd48605;
			16932: outdata = 32'd48604;
			16933: outdata = 32'd48603;
			16934: outdata = 32'd48602;
			16935: outdata = 32'd48601;
			16936: outdata = 32'd48600;
			16937: outdata = 32'd48599;
			16938: outdata = 32'd48598;
			16939: outdata = 32'd48597;
			16940: outdata = 32'd48596;
			16941: outdata = 32'd48595;
			16942: outdata = 32'd48594;
			16943: outdata = 32'd48593;
			16944: outdata = 32'd48592;
			16945: outdata = 32'd48591;
			16946: outdata = 32'd48590;
			16947: outdata = 32'd48589;
			16948: outdata = 32'd48588;
			16949: outdata = 32'd48587;
			16950: outdata = 32'd48586;
			16951: outdata = 32'd48585;
			16952: outdata = 32'd48584;
			16953: outdata = 32'd48583;
			16954: outdata = 32'd48582;
			16955: outdata = 32'd48581;
			16956: outdata = 32'd48580;
			16957: outdata = 32'd48579;
			16958: outdata = 32'd48578;
			16959: outdata = 32'd48577;
			16960: outdata = 32'd48576;
			16961: outdata = 32'd48575;
			16962: outdata = 32'd48574;
			16963: outdata = 32'd48573;
			16964: outdata = 32'd48572;
			16965: outdata = 32'd48571;
			16966: outdata = 32'd48570;
			16967: outdata = 32'd48569;
			16968: outdata = 32'd48568;
			16969: outdata = 32'd48567;
			16970: outdata = 32'd48566;
			16971: outdata = 32'd48565;
			16972: outdata = 32'd48564;
			16973: outdata = 32'd48563;
			16974: outdata = 32'd48562;
			16975: outdata = 32'd48561;
			16976: outdata = 32'd48560;
			16977: outdata = 32'd48559;
			16978: outdata = 32'd48558;
			16979: outdata = 32'd48557;
			16980: outdata = 32'd48556;
			16981: outdata = 32'd48555;
			16982: outdata = 32'd48554;
			16983: outdata = 32'd48553;
			16984: outdata = 32'd48552;
			16985: outdata = 32'd48551;
			16986: outdata = 32'd48550;
			16987: outdata = 32'd48549;
			16988: outdata = 32'd48548;
			16989: outdata = 32'd48547;
			16990: outdata = 32'd48546;
			16991: outdata = 32'd48545;
			16992: outdata = 32'd48544;
			16993: outdata = 32'd48543;
			16994: outdata = 32'd48542;
			16995: outdata = 32'd48541;
			16996: outdata = 32'd48540;
			16997: outdata = 32'd48539;
			16998: outdata = 32'd48538;
			16999: outdata = 32'd48537;
			17000: outdata = 32'd48536;
			17001: outdata = 32'd48535;
			17002: outdata = 32'd48534;
			17003: outdata = 32'd48533;
			17004: outdata = 32'd48532;
			17005: outdata = 32'd48531;
			17006: outdata = 32'd48530;
			17007: outdata = 32'd48529;
			17008: outdata = 32'd48528;
			17009: outdata = 32'd48527;
			17010: outdata = 32'd48526;
			17011: outdata = 32'd48525;
			17012: outdata = 32'd48524;
			17013: outdata = 32'd48523;
			17014: outdata = 32'd48522;
			17015: outdata = 32'd48521;
			17016: outdata = 32'd48520;
			17017: outdata = 32'd48519;
			17018: outdata = 32'd48518;
			17019: outdata = 32'd48517;
			17020: outdata = 32'd48516;
			17021: outdata = 32'd48515;
			17022: outdata = 32'd48514;
			17023: outdata = 32'd48513;
			17024: outdata = 32'd48512;
			17025: outdata = 32'd48511;
			17026: outdata = 32'd48510;
			17027: outdata = 32'd48509;
			17028: outdata = 32'd48508;
			17029: outdata = 32'd48507;
			17030: outdata = 32'd48506;
			17031: outdata = 32'd48505;
			17032: outdata = 32'd48504;
			17033: outdata = 32'd48503;
			17034: outdata = 32'd48502;
			17035: outdata = 32'd48501;
			17036: outdata = 32'd48500;
			17037: outdata = 32'd48499;
			17038: outdata = 32'd48498;
			17039: outdata = 32'd48497;
			17040: outdata = 32'd48496;
			17041: outdata = 32'd48495;
			17042: outdata = 32'd48494;
			17043: outdata = 32'd48493;
			17044: outdata = 32'd48492;
			17045: outdata = 32'd48491;
			17046: outdata = 32'd48490;
			17047: outdata = 32'd48489;
			17048: outdata = 32'd48488;
			17049: outdata = 32'd48487;
			17050: outdata = 32'd48486;
			17051: outdata = 32'd48485;
			17052: outdata = 32'd48484;
			17053: outdata = 32'd48483;
			17054: outdata = 32'd48482;
			17055: outdata = 32'd48481;
			17056: outdata = 32'd48480;
			17057: outdata = 32'd48479;
			17058: outdata = 32'd48478;
			17059: outdata = 32'd48477;
			17060: outdata = 32'd48476;
			17061: outdata = 32'd48475;
			17062: outdata = 32'd48474;
			17063: outdata = 32'd48473;
			17064: outdata = 32'd48472;
			17065: outdata = 32'd48471;
			17066: outdata = 32'd48470;
			17067: outdata = 32'd48469;
			17068: outdata = 32'd48468;
			17069: outdata = 32'd48467;
			17070: outdata = 32'd48466;
			17071: outdata = 32'd48465;
			17072: outdata = 32'd48464;
			17073: outdata = 32'd48463;
			17074: outdata = 32'd48462;
			17075: outdata = 32'd48461;
			17076: outdata = 32'd48460;
			17077: outdata = 32'd48459;
			17078: outdata = 32'd48458;
			17079: outdata = 32'd48457;
			17080: outdata = 32'd48456;
			17081: outdata = 32'd48455;
			17082: outdata = 32'd48454;
			17083: outdata = 32'd48453;
			17084: outdata = 32'd48452;
			17085: outdata = 32'd48451;
			17086: outdata = 32'd48450;
			17087: outdata = 32'd48449;
			17088: outdata = 32'd48448;
			17089: outdata = 32'd48447;
			17090: outdata = 32'd48446;
			17091: outdata = 32'd48445;
			17092: outdata = 32'd48444;
			17093: outdata = 32'd48443;
			17094: outdata = 32'd48442;
			17095: outdata = 32'd48441;
			17096: outdata = 32'd48440;
			17097: outdata = 32'd48439;
			17098: outdata = 32'd48438;
			17099: outdata = 32'd48437;
			17100: outdata = 32'd48436;
			17101: outdata = 32'd48435;
			17102: outdata = 32'd48434;
			17103: outdata = 32'd48433;
			17104: outdata = 32'd48432;
			17105: outdata = 32'd48431;
			17106: outdata = 32'd48430;
			17107: outdata = 32'd48429;
			17108: outdata = 32'd48428;
			17109: outdata = 32'd48427;
			17110: outdata = 32'd48426;
			17111: outdata = 32'd48425;
			17112: outdata = 32'd48424;
			17113: outdata = 32'd48423;
			17114: outdata = 32'd48422;
			17115: outdata = 32'd48421;
			17116: outdata = 32'd48420;
			17117: outdata = 32'd48419;
			17118: outdata = 32'd48418;
			17119: outdata = 32'd48417;
			17120: outdata = 32'd48416;
			17121: outdata = 32'd48415;
			17122: outdata = 32'd48414;
			17123: outdata = 32'd48413;
			17124: outdata = 32'd48412;
			17125: outdata = 32'd48411;
			17126: outdata = 32'd48410;
			17127: outdata = 32'd48409;
			17128: outdata = 32'd48408;
			17129: outdata = 32'd48407;
			17130: outdata = 32'd48406;
			17131: outdata = 32'd48405;
			17132: outdata = 32'd48404;
			17133: outdata = 32'd48403;
			17134: outdata = 32'd48402;
			17135: outdata = 32'd48401;
			17136: outdata = 32'd48400;
			17137: outdata = 32'd48399;
			17138: outdata = 32'd48398;
			17139: outdata = 32'd48397;
			17140: outdata = 32'd48396;
			17141: outdata = 32'd48395;
			17142: outdata = 32'd48394;
			17143: outdata = 32'd48393;
			17144: outdata = 32'd48392;
			17145: outdata = 32'd48391;
			17146: outdata = 32'd48390;
			17147: outdata = 32'd48389;
			17148: outdata = 32'd48388;
			17149: outdata = 32'd48387;
			17150: outdata = 32'd48386;
			17151: outdata = 32'd48385;
			17152: outdata = 32'd48384;
			17153: outdata = 32'd48383;
			17154: outdata = 32'd48382;
			17155: outdata = 32'd48381;
			17156: outdata = 32'd48380;
			17157: outdata = 32'd48379;
			17158: outdata = 32'd48378;
			17159: outdata = 32'd48377;
			17160: outdata = 32'd48376;
			17161: outdata = 32'd48375;
			17162: outdata = 32'd48374;
			17163: outdata = 32'd48373;
			17164: outdata = 32'd48372;
			17165: outdata = 32'd48371;
			17166: outdata = 32'd48370;
			17167: outdata = 32'd48369;
			17168: outdata = 32'd48368;
			17169: outdata = 32'd48367;
			17170: outdata = 32'd48366;
			17171: outdata = 32'd48365;
			17172: outdata = 32'd48364;
			17173: outdata = 32'd48363;
			17174: outdata = 32'd48362;
			17175: outdata = 32'd48361;
			17176: outdata = 32'd48360;
			17177: outdata = 32'd48359;
			17178: outdata = 32'd48358;
			17179: outdata = 32'd48357;
			17180: outdata = 32'd48356;
			17181: outdata = 32'd48355;
			17182: outdata = 32'd48354;
			17183: outdata = 32'd48353;
			17184: outdata = 32'd48352;
			17185: outdata = 32'd48351;
			17186: outdata = 32'd48350;
			17187: outdata = 32'd48349;
			17188: outdata = 32'd48348;
			17189: outdata = 32'd48347;
			17190: outdata = 32'd48346;
			17191: outdata = 32'd48345;
			17192: outdata = 32'd48344;
			17193: outdata = 32'd48343;
			17194: outdata = 32'd48342;
			17195: outdata = 32'd48341;
			17196: outdata = 32'd48340;
			17197: outdata = 32'd48339;
			17198: outdata = 32'd48338;
			17199: outdata = 32'd48337;
			17200: outdata = 32'd48336;
			17201: outdata = 32'd48335;
			17202: outdata = 32'd48334;
			17203: outdata = 32'd48333;
			17204: outdata = 32'd48332;
			17205: outdata = 32'd48331;
			17206: outdata = 32'd48330;
			17207: outdata = 32'd48329;
			17208: outdata = 32'd48328;
			17209: outdata = 32'd48327;
			17210: outdata = 32'd48326;
			17211: outdata = 32'd48325;
			17212: outdata = 32'd48324;
			17213: outdata = 32'd48323;
			17214: outdata = 32'd48322;
			17215: outdata = 32'd48321;
			17216: outdata = 32'd48320;
			17217: outdata = 32'd48319;
			17218: outdata = 32'd48318;
			17219: outdata = 32'd48317;
			17220: outdata = 32'd48316;
			17221: outdata = 32'd48315;
			17222: outdata = 32'd48314;
			17223: outdata = 32'd48313;
			17224: outdata = 32'd48312;
			17225: outdata = 32'd48311;
			17226: outdata = 32'd48310;
			17227: outdata = 32'd48309;
			17228: outdata = 32'd48308;
			17229: outdata = 32'd48307;
			17230: outdata = 32'd48306;
			17231: outdata = 32'd48305;
			17232: outdata = 32'd48304;
			17233: outdata = 32'd48303;
			17234: outdata = 32'd48302;
			17235: outdata = 32'd48301;
			17236: outdata = 32'd48300;
			17237: outdata = 32'd48299;
			17238: outdata = 32'd48298;
			17239: outdata = 32'd48297;
			17240: outdata = 32'd48296;
			17241: outdata = 32'd48295;
			17242: outdata = 32'd48294;
			17243: outdata = 32'd48293;
			17244: outdata = 32'd48292;
			17245: outdata = 32'd48291;
			17246: outdata = 32'd48290;
			17247: outdata = 32'd48289;
			17248: outdata = 32'd48288;
			17249: outdata = 32'd48287;
			17250: outdata = 32'd48286;
			17251: outdata = 32'd48285;
			17252: outdata = 32'd48284;
			17253: outdata = 32'd48283;
			17254: outdata = 32'd48282;
			17255: outdata = 32'd48281;
			17256: outdata = 32'd48280;
			17257: outdata = 32'd48279;
			17258: outdata = 32'd48278;
			17259: outdata = 32'd48277;
			17260: outdata = 32'd48276;
			17261: outdata = 32'd48275;
			17262: outdata = 32'd48274;
			17263: outdata = 32'd48273;
			17264: outdata = 32'd48272;
			17265: outdata = 32'd48271;
			17266: outdata = 32'd48270;
			17267: outdata = 32'd48269;
			17268: outdata = 32'd48268;
			17269: outdata = 32'd48267;
			17270: outdata = 32'd48266;
			17271: outdata = 32'd48265;
			17272: outdata = 32'd48264;
			17273: outdata = 32'd48263;
			17274: outdata = 32'd48262;
			17275: outdata = 32'd48261;
			17276: outdata = 32'd48260;
			17277: outdata = 32'd48259;
			17278: outdata = 32'd48258;
			17279: outdata = 32'd48257;
			17280: outdata = 32'd48256;
			17281: outdata = 32'd48255;
			17282: outdata = 32'd48254;
			17283: outdata = 32'd48253;
			17284: outdata = 32'd48252;
			17285: outdata = 32'd48251;
			17286: outdata = 32'd48250;
			17287: outdata = 32'd48249;
			17288: outdata = 32'd48248;
			17289: outdata = 32'd48247;
			17290: outdata = 32'd48246;
			17291: outdata = 32'd48245;
			17292: outdata = 32'd48244;
			17293: outdata = 32'd48243;
			17294: outdata = 32'd48242;
			17295: outdata = 32'd48241;
			17296: outdata = 32'd48240;
			17297: outdata = 32'd48239;
			17298: outdata = 32'd48238;
			17299: outdata = 32'd48237;
			17300: outdata = 32'd48236;
			17301: outdata = 32'd48235;
			17302: outdata = 32'd48234;
			17303: outdata = 32'd48233;
			17304: outdata = 32'd48232;
			17305: outdata = 32'd48231;
			17306: outdata = 32'd48230;
			17307: outdata = 32'd48229;
			17308: outdata = 32'd48228;
			17309: outdata = 32'd48227;
			17310: outdata = 32'd48226;
			17311: outdata = 32'd48225;
			17312: outdata = 32'd48224;
			17313: outdata = 32'd48223;
			17314: outdata = 32'd48222;
			17315: outdata = 32'd48221;
			17316: outdata = 32'd48220;
			17317: outdata = 32'd48219;
			17318: outdata = 32'd48218;
			17319: outdata = 32'd48217;
			17320: outdata = 32'd48216;
			17321: outdata = 32'd48215;
			17322: outdata = 32'd48214;
			17323: outdata = 32'd48213;
			17324: outdata = 32'd48212;
			17325: outdata = 32'd48211;
			17326: outdata = 32'd48210;
			17327: outdata = 32'd48209;
			17328: outdata = 32'd48208;
			17329: outdata = 32'd48207;
			17330: outdata = 32'd48206;
			17331: outdata = 32'd48205;
			17332: outdata = 32'd48204;
			17333: outdata = 32'd48203;
			17334: outdata = 32'd48202;
			17335: outdata = 32'd48201;
			17336: outdata = 32'd48200;
			17337: outdata = 32'd48199;
			17338: outdata = 32'd48198;
			17339: outdata = 32'd48197;
			17340: outdata = 32'd48196;
			17341: outdata = 32'd48195;
			17342: outdata = 32'd48194;
			17343: outdata = 32'd48193;
			17344: outdata = 32'd48192;
			17345: outdata = 32'd48191;
			17346: outdata = 32'd48190;
			17347: outdata = 32'd48189;
			17348: outdata = 32'd48188;
			17349: outdata = 32'd48187;
			17350: outdata = 32'd48186;
			17351: outdata = 32'd48185;
			17352: outdata = 32'd48184;
			17353: outdata = 32'd48183;
			17354: outdata = 32'd48182;
			17355: outdata = 32'd48181;
			17356: outdata = 32'd48180;
			17357: outdata = 32'd48179;
			17358: outdata = 32'd48178;
			17359: outdata = 32'd48177;
			17360: outdata = 32'd48176;
			17361: outdata = 32'd48175;
			17362: outdata = 32'd48174;
			17363: outdata = 32'd48173;
			17364: outdata = 32'd48172;
			17365: outdata = 32'd48171;
			17366: outdata = 32'd48170;
			17367: outdata = 32'd48169;
			17368: outdata = 32'd48168;
			17369: outdata = 32'd48167;
			17370: outdata = 32'd48166;
			17371: outdata = 32'd48165;
			17372: outdata = 32'd48164;
			17373: outdata = 32'd48163;
			17374: outdata = 32'd48162;
			17375: outdata = 32'd48161;
			17376: outdata = 32'd48160;
			17377: outdata = 32'd48159;
			17378: outdata = 32'd48158;
			17379: outdata = 32'd48157;
			17380: outdata = 32'd48156;
			17381: outdata = 32'd48155;
			17382: outdata = 32'd48154;
			17383: outdata = 32'd48153;
			17384: outdata = 32'd48152;
			17385: outdata = 32'd48151;
			17386: outdata = 32'd48150;
			17387: outdata = 32'd48149;
			17388: outdata = 32'd48148;
			17389: outdata = 32'd48147;
			17390: outdata = 32'd48146;
			17391: outdata = 32'd48145;
			17392: outdata = 32'd48144;
			17393: outdata = 32'd48143;
			17394: outdata = 32'd48142;
			17395: outdata = 32'd48141;
			17396: outdata = 32'd48140;
			17397: outdata = 32'd48139;
			17398: outdata = 32'd48138;
			17399: outdata = 32'd48137;
			17400: outdata = 32'd48136;
			17401: outdata = 32'd48135;
			17402: outdata = 32'd48134;
			17403: outdata = 32'd48133;
			17404: outdata = 32'd48132;
			17405: outdata = 32'd48131;
			17406: outdata = 32'd48130;
			17407: outdata = 32'd48129;
			17408: outdata = 32'd48128;
			17409: outdata = 32'd48127;
			17410: outdata = 32'd48126;
			17411: outdata = 32'd48125;
			17412: outdata = 32'd48124;
			17413: outdata = 32'd48123;
			17414: outdata = 32'd48122;
			17415: outdata = 32'd48121;
			17416: outdata = 32'd48120;
			17417: outdata = 32'd48119;
			17418: outdata = 32'd48118;
			17419: outdata = 32'd48117;
			17420: outdata = 32'd48116;
			17421: outdata = 32'd48115;
			17422: outdata = 32'd48114;
			17423: outdata = 32'd48113;
			17424: outdata = 32'd48112;
			17425: outdata = 32'd48111;
			17426: outdata = 32'd48110;
			17427: outdata = 32'd48109;
			17428: outdata = 32'd48108;
			17429: outdata = 32'd48107;
			17430: outdata = 32'd48106;
			17431: outdata = 32'd48105;
			17432: outdata = 32'd48104;
			17433: outdata = 32'd48103;
			17434: outdata = 32'd48102;
			17435: outdata = 32'd48101;
			17436: outdata = 32'd48100;
			17437: outdata = 32'd48099;
			17438: outdata = 32'd48098;
			17439: outdata = 32'd48097;
			17440: outdata = 32'd48096;
			17441: outdata = 32'd48095;
			17442: outdata = 32'd48094;
			17443: outdata = 32'd48093;
			17444: outdata = 32'd48092;
			17445: outdata = 32'd48091;
			17446: outdata = 32'd48090;
			17447: outdata = 32'd48089;
			17448: outdata = 32'd48088;
			17449: outdata = 32'd48087;
			17450: outdata = 32'd48086;
			17451: outdata = 32'd48085;
			17452: outdata = 32'd48084;
			17453: outdata = 32'd48083;
			17454: outdata = 32'd48082;
			17455: outdata = 32'd48081;
			17456: outdata = 32'd48080;
			17457: outdata = 32'd48079;
			17458: outdata = 32'd48078;
			17459: outdata = 32'd48077;
			17460: outdata = 32'd48076;
			17461: outdata = 32'd48075;
			17462: outdata = 32'd48074;
			17463: outdata = 32'd48073;
			17464: outdata = 32'd48072;
			17465: outdata = 32'd48071;
			17466: outdata = 32'd48070;
			17467: outdata = 32'd48069;
			17468: outdata = 32'd48068;
			17469: outdata = 32'd48067;
			17470: outdata = 32'd48066;
			17471: outdata = 32'd48065;
			17472: outdata = 32'd48064;
			17473: outdata = 32'd48063;
			17474: outdata = 32'd48062;
			17475: outdata = 32'd48061;
			17476: outdata = 32'd48060;
			17477: outdata = 32'd48059;
			17478: outdata = 32'd48058;
			17479: outdata = 32'd48057;
			17480: outdata = 32'd48056;
			17481: outdata = 32'd48055;
			17482: outdata = 32'd48054;
			17483: outdata = 32'd48053;
			17484: outdata = 32'd48052;
			17485: outdata = 32'd48051;
			17486: outdata = 32'd48050;
			17487: outdata = 32'd48049;
			17488: outdata = 32'd48048;
			17489: outdata = 32'd48047;
			17490: outdata = 32'd48046;
			17491: outdata = 32'd48045;
			17492: outdata = 32'd48044;
			17493: outdata = 32'd48043;
			17494: outdata = 32'd48042;
			17495: outdata = 32'd48041;
			17496: outdata = 32'd48040;
			17497: outdata = 32'd48039;
			17498: outdata = 32'd48038;
			17499: outdata = 32'd48037;
			17500: outdata = 32'd48036;
			17501: outdata = 32'd48035;
			17502: outdata = 32'd48034;
			17503: outdata = 32'd48033;
			17504: outdata = 32'd48032;
			17505: outdata = 32'd48031;
			17506: outdata = 32'd48030;
			17507: outdata = 32'd48029;
			17508: outdata = 32'd48028;
			17509: outdata = 32'd48027;
			17510: outdata = 32'd48026;
			17511: outdata = 32'd48025;
			17512: outdata = 32'd48024;
			17513: outdata = 32'd48023;
			17514: outdata = 32'd48022;
			17515: outdata = 32'd48021;
			17516: outdata = 32'd48020;
			17517: outdata = 32'd48019;
			17518: outdata = 32'd48018;
			17519: outdata = 32'd48017;
			17520: outdata = 32'd48016;
			17521: outdata = 32'd48015;
			17522: outdata = 32'd48014;
			17523: outdata = 32'd48013;
			17524: outdata = 32'd48012;
			17525: outdata = 32'd48011;
			17526: outdata = 32'd48010;
			17527: outdata = 32'd48009;
			17528: outdata = 32'd48008;
			17529: outdata = 32'd48007;
			17530: outdata = 32'd48006;
			17531: outdata = 32'd48005;
			17532: outdata = 32'd48004;
			17533: outdata = 32'd48003;
			17534: outdata = 32'd48002;
			17535: outdata = 32'd48001;
			17536: outdata = 32'd48000;
			17537: outdata = 32'd47999;
			17538: outdata = 32'd47998;
			17539: outdata = 32'd47997;
			17540: outdata = 32'd47996;
			17541: outdata = 32'd47995;
			17542: outdata = 32'd47994;
			17543: outdata = 32'd47993;
			17544: outdata = 32'd47992;
			17545: outdata = 32'd47991;
			17546: outdata = 32'd47990;
			17547: outdata = 32'd47989;
			17548: outdata = 32'd47988;
			17549: outdata = 32'd47987;
			17550: outdata = 32'd47986;
			17551: outdata = 32'd47985;
			17552: outdata = 32'd47984;
			17553: outdata = 32'd47983;
			17554: outdata = 32'd47982;
			17555: outdata = 32'd47981;
			17556: outdata = 32'd47980;
			17557: outdata = 32'd47979;
			17558: outdata = 32'd47978;
			17559: outdata = 32'd47977;
			17560: outdata = 32'd47976;
			17561: outdata = 32'd47975;
			17562: outdata = 32'd47974;
			17563: outdata = 32'd47973;
			17564: outdata = 32'd47972;
			17565: outdata = 32'd47971;
			17566: outdata = 32'd47970;
			17567: outdata = 32'd47969;
			17568: outdata = 32'd47968;
			17569: outdata = 32'd47967;
			17570: outdata = 32'd47966;
			17571: outdata = 32'd47965;
			17572: outdata = 32'd47964;
			17573: outdata = 32'd47963;
			17574: outdata = 32'd47962;
			17575: outdata = 32'd47961;
			17576: outdata = 32'd47960;
			17577: outdata = 32'd47959;
			17578: outdata = 32'd47958;
			17579: outdata = 32'd47957;
			17580: outdata = 32'd47956;
			17581: outdata = 32'd47955;
			17582: outdata = 32'd47954;
			17583: outdata = 32'd47953;
			17584: outdata = 32'd47952;
			17585: outdata = 32'd47951;
			17586: outdata = 32'd47950;
			17587: outdata = 32'd47949;
			17588: outdata = 32'd47948;
			17589: outdata = 32'd47947;
			17590: outdata = 32'd47946;
			17591: outdata = 32'd47945;
			17592: outdata = 32'd47944;
			17593: outdata = 32'd47943;
			17594: outdata = 32'd47942;
			17595: outdata = 32'd47941;
			17596: outdata = 32'd47940;
			17597: outdata = 32'd47939;
			17598: outdata = 32'd47938;
			17599: outdata = 32'd47937;
			17600: outdata = 32'd47936;
			17601: outdata = 32'd47935;
			17602: outdata = 32'd47934;
			17603: outdata = 32'd47933;
			17604: outdata = 32'd47932;
			17605: outdata = 32'd47931;
			17606: outdata = 32'd47930;
			17607: outdata = 32'd47929;
			17608: outdata = 32'd47928;
			17609: outdata = 32'd47927;
			17610: outdata = 32'd47926;
			17611: outdata = 32'd47925;
			17612: outdata = 32'd47924;
			17613: outdata = 32'd47923;
			17614: outdata = 32'd47922;
			17615: outdata = 32'd47921;
			17616: outdata = 32'd47920;
			17617: outdata = 32'd47919;
			17618: outdata = 32'd47918;
			17619: outdata = 32'd47917;
			17620: outdata = 32'd47916;
			17621: outdata = 32'd47915;
			17622: outdata = 32'd47914;
			17623: outdata = 32'd47913;
			17624: outdata = 32'd47912;
			17625: outdata = 32'd47911;
			17626: outdata = 32'd47910;
			17627: outdata = 32'd47909;
			17628: outdata = 32'd47908;
			17629: outdata = 32'd47907;
			17630: outdata = 32'd47906;
			17631: outdata = 32'd47905;
			17632: outdata = 32'd47904;
			17633: outdata = 32'd47903;
			17634: outdata = 32'd47902;
			17635: outdata = 32'd47901;
			17636: outdata = 32'd47900;
			17637: outdata = 32'd47899;
			17638: outdata = 32'd47898;
			17639: outdata = 32'd47897;
			17640: outdata = 32'd47896;
			17641: outdata = 32'd47895;
			17642: outdata = 32'd47894;
			17643: outdata = 32'd47893;
			17644: outdata = 32'd47892;
			17645: outdata = 32'd47891;
			17646: outdata = 32'd47890;
			17647: outdata = 32'd47889;
			17648: outdata = 32'd47888;
			17649: outdata = 32'd47887;
			17650: outdata = 32'd47886;
			17651: outdata = 32'd47885;
			17652: outdata = 32'd47884;
			17653: outdata = 32'd47883;
			17654: outdata = 32'd47882;
			17655: outdata = 32'd47881;
			17656: outdata = 32'd47880;
			17657: outdata = 32'd47879;
			17658: outdata = 32'd47878;
			17659: outdata = 32'd47877;
			17660: outdata = 32'd47876;
			17661: outdata = 32'd47875;
			17662: outdata = 32'd47874;
			17663: outdata = 32'd47873;
			17664: outdata = 32'd47872;
			17665: outdata = 32'd47871;
			17666: outdata = 32'd47870;
			17667: outdata = 32'd47869;
			17668: outdata = 32'd47868;
			17669: outdata = 32'd47867;
			17670: outdata = 32'd47866;
			17671: outdata = 32'd47865;
			17672: outdata = 32'd47864;
			17673: outdata = 32'd47863;
			17674: outdata = 32'd47862;
			17675: outdata = 32'd47861;
			17676: outdata = 32'd47860;
			17677: outdata = 32'd47859;
			17678: outdata = 32'd47858;
			17679: outdata = 32'd47857;
			17680: outdata = 32'd47856;
			17681: outdata = 32'd47855;
			17682: outdata = 32'd47854;
			17683: outdata = 32'd47853;
			17684: outdata = 32'd47852;
			17685: outdata = 32'd47851;
			17686: outdata = 32'd47850;
			17687: outdata = 32'd47849;
			17688: outdata = 32'd47848;
			17689: outdata = 32'd47847;
			17690: outdata = 32'd47846;
			17691: outdata = 32'd47845;
			17692: outdata = 32'd47844;
			17693: outdata = 32'd47843;
			17694: outdata = 32'd47842;
			17695: outdata = 32'd47841;
			17696: outdata = 32'd47840;
			17697: outdata = 32'd47839;
			17698: outdata = 32'd47838;
			17699: outdata = 32'd47837;
			17700: outdata = 32'd47836;
			17701: outdata = 32'd47835;
			17702: outdata = 32'd47834;
			17703: outdata = 32'd47833;
			17704: outdata = 32'd47832;
			17705: outdata = 32'd47831;
			17706: outdata = 32'd47830;
			17707: outdata = 32'd47829;
			17708: outdata = 32'd47828;
			17709: outdata = 32'd47827;
			17710: outdata = 32'd47826;
			17711: outdata = 32'd47825;
			17712: outdata = 32'd47824;
			17713: outdata = 32'd47823;
			17714: outdata = 32'd47822;
			17715: outdata = 32'd47821;
			17716: outdata = 32'd47820;
			17717: outdata = 32'd47819;
			17718: outdata = 32'd47818;
			17719: outdata = 32'd47817;
			17720: outdata = 32'd47816;
			17721: outdata = 32'd47815;
			17722: outdata = 32'd47814;
			17723: outdata = 32'd47813;
			17724: outdata = 32'd47812;
			17725: outdata = 32'd47811;
			17726: outdata = 32'd47810;
			17727: outdata = 32'd47809;
			17728: outdata = 32'd47808;
			17729: outdata = 32'd47807;
			17730: outdata = 32'd47806;
			17731: outdata = 32'd47805;
			17732: outdata = 32'd47804;
			17733: outdata = 32'd47803;
			17734: outdata = 32'd47802;
			17735: outdata = 32'd47801;
			17736: outdata = 32'd47800;
			17737: outdata = 32'd47799;
			17738: outdata = 32'd47798;
			17739: outdata = 32'd47797;
			17740: outdata = 32'd47796;
			17741: outdata = 32'd47795;
			17742: outdata = 32'd47794;
			17743: outdata = 32'd47793;
			17744: outdata = 32'd47792;
			17745: outdata = 32'd47791;
			17746: outdata = 32'd47790;
			17747: outdata = 32'd47789;
			17748: outdata = 32'd47788;
			17749: outdata = 32'd47787;
			17750: outdata = 32'd47786;
			17751: outdata = 32'd47785;
			17752: outdata = 32'd47784;
			17753: outdata = 32'd47783;
			17754: outdata = 32'd47782;
			17755: outdata = 32'd47781;
			17756: outdata = 32'd47780;
			17757: outdata = 32'd47779;
			17758: outdata = 32'd47778;
			17759: outdata = 32'd47777;
			17760: outdata = 32'd47776;
			17761: outdata = 32'd47775;
			17762: outdata = 32'd47774;
			17763: outdata = 32'd47773;
			17764: outdata = 32'd47772;
			17765: outdata = 32'd47771;
			17766: outdata = 32'd47770;
			17767: outdata = 32'd47769;
			17768: outdata = 32'd47768;
			17769: outdata = 32'd47767;
			17770: outdata = 32'd47766;
			17771: outdata = 32'd47765;
			17772: outdata = 32'd47764;
			17773: outdata = 32'd47763;
			17774: outdata = 32'd47762;
			17775: outdata = 32'd47761;
			17776: outdata = 32'd47760;
			17777: outdata = 32'd47759;
			17778: outdata = 32'd47758;
			17779: outdata = 32'd47757;
			17780: outdata = 32'd47756;
			17781: outdata = 32'd47755;
			17782: outdata = 32'd47754;
			17783: outdata = 32'd47753;
			17784: outdata = 32'd47752;
			17785: outdata = 32'd47751;
			17786: outdata = 32'd47750;
			17787: outdata = 32'd47749;
			17788: outdata = 32'd47748;
			17789: outdata = 32'd47747;
			17790: outdata = 32'd47746;
			17791: outdata = 32'd47745;
			17792: outdata = 32'd47744;
			17793: outdata = 32'd47743;
			17794: outdata = 32'd47742;
			17795: outdata = 32'd47741;
			17796: outdata = 32'd47740;
			17797: outdata = 32'd47739;
			17798: outdata = 32'd47738;
			17799: outdata = 32'd47737;
			17800: outdata = 32'd47736;
			17801: outdata = 32'd47735;
			17802: outdata = 32'd47734;
			17803: outdata = 32'd47733;
			17804: outdata = 32'd47732;
			17805: outdata = 32'd47731;
			17806: outdata = 32'd47730;
			17807: outdata = 32'd47729;
			17808: outdata = 32'd47728;
			17809: outdata = 32'd47727;
			17810: outdata = 32'd47726;
			17811: outdata = 32'd47725;
			17812: outdata = 32'd47724;
			17813: outdata = 32'd47723;
			17814: outdata = 32'd47722;
			17815: outdata = 32'd47721;
			17816: outdata = 32'd47720;
			17817: outdata = 32'd47719;
			17818: outdata = 32'd47718;
			17819: outdata = 32'd47717;
			17820: outdata = 32'd47716;
			17821: outdata = 32'd47715;
			17822: outdata = 32'd47714;
			17823: outdata = 32'd47713;
			17824: outdata = 32'd47712;
			17825: outdata = 32'd47711;
			17826: outdata = 32'd47710;
			17827: outdata = 32'd47709;
			17828: outdata = 32'd47708;
			17829: outdata = 32'd47707;
			17830: outdata = 32'd47706;
			17831: outdata = 32'd47705;
			17832: outdata = 32'd47704;
			17833: outdata = 32'd47703;
			17834: outdata = 32'd47702;
			17835: outdata = 32'd47701;
			17836: outdata = 32'd47700;
			17837: outdata = 32'd47699;
			17838: outdata = 32'd47698;
			17839: outdata = 32'd47697;
			17840: outdata = 32'd47696;
			17841: outdata = 32'd47695;
			17842: outdata = 32'd47694;
			17843: outdata = 32'd47693;
			17844: outdata = 32'd47692;
			17845: outdata = 32'd47691;
			17846: outdata = 32'd47690;
			17847: outdata = 32'd47689;
			17848: outdata = 32'd47688;
			17849: outdata = 32'd47687;
			17850: outdata = 32'd47686;
			17851: outdata = 32'd47685;
			17852: outdata = 32'd47684;
			17853: outdata = 32'd47683;
			17854: outdata = 32'd47682;
			17855: outdata = 32'd47681;
			17856: outdata = 32'd47680;
			17857: outdata = 32'd47679;
			17858: outdata = 32'd47678;
			17859: outdata = 32'd47677;
			17860: outdata = 32'd47676;
			17861: outdata = 32'd47675;
			17862: outdata = 32'd47674;
			17863: outdata = 32'd47673;
			17864: outdata = 32'd47672;
			17865: outdata = 32'd47671;
			17866: outdata = 32'd47670;
			17867: outdata = 32'd47669;
			17868: outdata = 32'd47668;
			17869: outdata = 32'd47667;
			17870: outdata = 32'd47666;
			17871: outdata = 32'd47665;
			17872: outdata = 32'd47664;
			17873: outdata = 32'd47663;
			17874: outdata = 32'd47662;
			17875: outdata = 32'd47661;
			17876: outdata = 32'd47660;
			17877: outdata = 32'd47659;
			17878: outdata = 32'd47658;
			17879: outdata = 32'd47657;
			17880: outdata = 32'd47656;
			17881: outdata = 32'd47655;
			17882: outdata = 32'd47654;
			17883: outdata = 32'd47653;
			17884: outdata = 32'd47652;
			17885: outdata = 32'd47651;
			17886: outdata = 32'd47650;
			17887: outdata = 32'd47649;
			17888: outdata = 32'd47648;
			17889: outdata = 32'd47647;
			17890: outdata = 32'd47646;
			17891: outdata = 32'd47645;
			17892: outdata = 32'd47644;
			17893: outdata = 32'd47643;
			17894: outdata = 32'd47642;
			17895: outdata = 32'd47641;
			17896: outdata = 32'd47640;
			17897: outdata = 32'd47639;
			17898: outdata = 32'd47638;
			17899: outdata = 32'd47637;
			17900: outdata = 32'd47636;
			17901: outdata = 32'd47635;
			17902: outdata = 32'd47634;
			17903: outdata = 32'd47633;
			17904: outdata = 32'd47632;
			17905: outdata = 32'd47631;
			17906: outdata = 32'd47630;
			17907: outdata = 32'd47629;
			17908: outdata = 32'd47628;
			17909: outdata = 32'd47627;
			17910: outdata = 32'd47626;
			17911: outdata = 32'd47625;
			17912: outdata = 32'd47624;
			17913: outdata = 32'd47623;
			17914: outdata = 32'd47622;
			17915: outdata = 32'd47621;
			17916: outdata = 32'd47620;
			17917: outdata = 32'd47619;
			17918: outdata = 32'd47618;
			17919: outdata = 32'd47617;
			17920: outdata = 32'd47616;
			17921: outdata = 32'd47615;
			17922: outdata = 32'd47614;
			17923: outdata = 32'd47613;
			17924: outdata = 32'd47612;
			17925: outdata = 32'd47611;
			17926: outdata = 32'd47610;
			17927: outdata = 32'd47609;
			17928: outdata = 32'd47608;
			17929: outdata = 32'd47607;
			17930: outdata = 32'd47606;
			17931: outdata = 32'd47605;
			17932: outdata = 32'd47604;
			17933: outdata = 32'd47603;
			17934: outdata = 32'd47602;
			17935: outdata = 32'd47601;
			17936: outdata = 32'd47600;
			17937: outdata = 32'd47599;
			17938: outdata = 32'd47598;
			17939: outdata = 32'd47597;
			17940: outdata = 32'd47596;
			17941: outdata = 32'd47595;
			17942: outdata = 32'd47594;
			17943: outdata = 32'd47593;
			17944: outdata = 32'd47592;
			17945: outdata = 32'd47591;
			17946: outdata = 32'd47590;
			17947: outdata = 32'd47589;
			17948: outdata = 32'd47588;
			17949: outdata = 32'd47587;
			17950: outdata = 32'd47586;
			17951: outdata = 32'd47585;
			17952: outdata = 32'd47584;
			17953: outdata = 32'd47583;
			17954: outdata = 32'd47582;
			17955: outdata = 32'd47581;
			17956: outdata = 32'd47580;
			17957: outdata = 32'd47579;
			17958: outdata = 32'd47578;
			17959: outdata = 32'd47577;
			17960: outdata = 32'd47576;
			17961: outdata = 32'd47575;
			17962: outdata = 32'd47574;
			17963: outdata = 32'd47573;
			17964: outdata = 32'd47572;
			17965: outdata = 32'd47571;
			17966: outdata = 32'd47570;
			17967: outdata = 32'd47569;
			17968: outdata = 32'd47568;
			17969: outdata = 32'd47567;
			17970: outdata = 32'd47566;
			17971: outdata = 32'd47565;
			17972: outdata = 32'd47564;
			17973: outdata = 32'd47563;
			17974: outdata = 32'd47562;
			17975: outdata = 32'd47561;
			17976: outdata = 32'd47560;
			17977: outdata = 32'd47559;
			17978: outdata = 32'd47558;
			17979: outdata = 32'd47557;
			17980: outdata = 32'd47556;
			17981: outdata = 32'd47555;
			17982: outdata = 32'd47554;
			17983: outdata = 32'd47553;
			17984: outdata = 32'd47552;
			17985: outdata = 32'd47551;
			17986: outdata = 32'd47550;
			17987: outdata = 32'd47549;
			17988: outdata = 32'd47548;
			17989: outdata = 32'd47547;
			17990: outdata = 32'd47546;
			17991: outdata = 32'd47545;
			17992: outdata = 32'd47544;
			17993: outdata = 32'd47543;
			17994: outdata = 32'd47542;
			17995: outdata = 32'd47541;
			17996: outdata = 32'd47540;
			17997: outdata = 32'd47539;
			17998: outdata = 32'd47538;
			17999: outdata = 32'd47537;
			18000: outdata = 32'd47536;
			18001: outdata = 32'd47535;
			18002: outdata = 32'd47534;
			18003: outdata = 32'd47533;
			18004: outdata = 32'd47532;
			18005: outdata = 32'd47531;
			18006: outdata = 32'd47530;
			18007: outdata = 32'd47529;
			18008: outdata = 32'd47528;
			18009: outdata = 32'd47527;
			18010: outdata = 32'd47526;
			18011: outdata = 32'd47525;
			18012: outdata = 32'd47524;
			18013: outdata = 32'd47523;
			18014: outdata = 32'd47522;
			18015: outdata = 32'd47521;
			18016: outdata = 32'd47520;
			18017: outdata = 32'd47519;
			18018: outdata = 32'd47518;
			18019: outdata = 32'd47517;
			18020: outdata = 32'd47516;
			18021: outdata = 32'd47515;
			18022: outdata = 32'd47514;
			18023: outdata = 32'd47513;
			18024: outdata = 32'd47512;
			18025: outdata = 32'd47511;
			18026: outdata = 32'd47510;
			18027: outdata = 32'd47509;
			18028: outdata = 32'd47508;
			18029: outdata = 32'd47507;
			18030: outdata = 32'd47506;
			18031: outdata = 32'd47505;
			18032: outdata = 32'd47504;
			18033: outdata = 32'd47503;
			18034: outdata = 32'd47502;
			18035: outdata = 32'd47501;
			18036: outdata = 32'd47500;
			18037: outdata = 32'd47499;
			18038: outdata = 32'd47498;
			18039: outdata = 32'd47497;
			18040: outdata = 32'd47496;
			18041: outdata = 32'd47495;
			18042: outdata = 32'd47494;
			18043: outdata = 32'd47493;
			18044: outdata = 32'd47492;
			18045: outdata = 32'd47491;
			18046: outdata = 32'd47490;
			18047: outdata = 32'd47489;
			18048: outdata = 32'd47488;
			18049: outdata = 32'd47487;
			18050: outdata = 32'd47486;
			18051: outdata = 32'd47485;
			18052: outdata = 32'd47484;
			18053: outdata = 32'd47483;
			18054: outdata = 32'd47482;
			18055: outdata = 32'd47481;
			18056: outdata = 32'd47480;
			18057: outdata = 32'd47479;
			18058: outdata = 32'd47478;
			18059: outdata = 32'd47477;
			18060: outdata = 32'd47476;
			18061: outdata = 32'd47475;
			18062: outdata = 32'd47474;
			18063: outdata = 32'd47473;
			18064: outdata = 32'd47472;
			18065: outdata = 32'd47471;
			18066: outdata = 32'd47470;
			18067: outdata = 32'd47469;
			18068: outdata = 32'd47468;
			18069: outdata = 32'd47467;
			18070: outdata = 32'd47466;
			18071: outdata = 32'd47465;
			18072: outdata = 32'd47464;
			18073: outdata = 32'd47463;
			18074: outdata = 32'd47462;
			18075: outdata = 32'd47461;
			18076: outdata = 32'd47460;
			18077: outdata = 32'd47459;
			18078: outdata = 32'd47458;
			18079: outdata = 32'd47457;
			18080: outdata = 32'd47456;
			18081: outdata = 32'd47455;
			18082: outdata = 32'd47454;
			18083: outdata = 32'd47453;
			18084: outdata = 32'd47452;
			18085: outdata = 32'd47451;
			18086: outdata = 32'd47450;
			18087: outdata = 32'd47449;
			18088: outdata = 32'd47448;
			18089: outdata = 32'd47447;
			18090: outdata = 32'd47446;
			18091: outdata = 32'd47445;
			18092: outdata = 32'd47444;
			18093: outdata = 32'd47443;
			18094: outdata = 32'd47442;
			18095: outdata = 32'd47441;
			18096: outdata = 32'd47440;
			18097: outdata = 32'd47439;
			18098: outdata = 32'd47438;
			18099: outdata = 32'd47437;
			18100: outdata = 32'd47436;
			18101: outdata = 32'd47435;
			18102: outdata = 32'd47434;
			18103: outdata = 32'd47433;
			18104: outdata = 32'd47432;
			18105: outdata = 32'd47431;
			18106: outdata = 32'd47430;
			18107: outdata = 32'd47429;
			18108: outdata = 32'd47428;
			18109: outdata = 32'd47427;
			18110: outdata = 32'd47426;
			18111: outdata = 32'd47425;
			18112: outdata = 32'd47424;
			18113: outdata = 32'd47423;
			18114: outdata = 32'd47422;
			18115: outdata = 32'd47421;
			18116: outdata = 32'd47420;
			18117: outdata = 32'd47419;
			18118: outdata = 32'd47418;
			18119: outdata = 32'd47417;
			18120: outdata = 32'd47416;
			18121: outdata = 32'd47415;
			18122: outdata = 32'd47414;
			18123: outdata = 32'd47413;
			18124: outdata = 32'd47412;
			18125: outdata = 32'd47411;
			18126: outdata = 32'd47410;
			18127: outdata = 32'd47409;
			18128: outdata = 32'd47408;
			18129: outdata = 32'd47407;
			18130: outdata = 32'd47406;
			18131: outdata = 32'd47405;
			18132: outdata = 32'd47404;
			18133: outdata = 32'd47403;
			18134: outdata = 32'd47402;
			18135: outdata = 32'd47401;
			18136: outdata = 32'd47400;
			18137: outdata = 32'd47399;
			18138: outdata = 32'd47398;
			18139: outdata = 32'd47397;
			18140: outdata = 32'd47396;
			18141: outdata = 32'd47395;
			18142: outdata = 32'd47394;
			18143: outdata = 32'd47393;
			18144: outdata = 32'd47392;
			18145: outdata = 32'd47391;
			18146: outdata = 32'd47390;
			18147: outdata = 32'd47389;
			18148: outdata = 32'd47388;
			18149: outdata = 32'd47387;
			18150: outdata = 32'd47386;
			18151: outdata = 32'd47385;
			18152: outdata = 32'd47384;
			18153: outdata = 32'd47383;
			18154: outdata = 32'd47382;
			18155: outdata = 32'd47381;
			18156: outdata = 32'd47380;
			18157: outdata = 32'd47379;
			18158: outdata = 32'd47378;
			18159: outdata = 32'd47377;
			18160: outdata = 32'd47376;
			18161: outdata = 32'd47375;
			18162: outdata = 32'd47374;
			18163: outdata = 32'd47373;
			18164: outdata = 32'd47372;
			18165: outdata = 32'd47371;
			18166: outdata = 32'd47370;
			18167: outdata = 32'd47369;
			18168: outdata = 32'd47368;
			18169: outdata = 32'd47367;
			18170: outdata = 32'd47366;
			18171: outdata = 32'd47365;
			18172: outdata = 32'd47364;
			18173: outdata = 32'd47363;
			18174: outdata = 32'd47362;
			18175: outdata = 32'd47361;
			18176: outdata = 32'd47360;
			18177: outdata = 32'd47359;
			18178: outdata = 32'd47358;
			18179: outdata = 32'd47357;
			18180: outdata = 32'd47356;
			18181: outdata = 32'd47355;
			18182: outdata = 32'd47354;
			18183: outdata = 32'd47353;
			18184: outdata = 32'd47352;
			18185: outdata = 32'd47351;
			18186: outdata = 32'd47350;
			18187: outdata = 32'd47349;
			18188: outdata = 32'd47348;
			18189: outdata = 32'd47347;
			18190: outdata = 32'd47346;
			18191: outdata = 32'd47345;
			18192: outdata = 32'd47344;
			18193: outdata = 32'd47343;
			18194: outdata = 32'd47342;
			18195: outdata = 32'd47341;
			18196: outdata = 32'd47340;
			18197: outdata = 32'd47339;
			18198: outdata = 32'd47338;
			18199: outdata = 32'd47337;
			18200: outdata = 32'd47336;
			18201: outdata = 32'd47335;
			18202: outdata = 32'd47334;
			18203: outdata = 32'd47333;
			18204: outdata = 32'd47332;
			18205: outdata = 32'd47331;
			18206: outdata = 32'd47330;
			18207: outdata = 32'd47329;
			18208: outdata = 32'd47328;
			18209: outdata = 32'd47327;
			18210: outdata = 32'd47326;
			18211: outdata = 32'd47325;
			18212: outdata = 32'd47324;
			18213: outdata = 32'd47323;
			18214: outdata = 32'd47322;
			18215: outdata = 32'd47321;
			18216: outdata = 32'd47320;
			18217: outdata = 32'd47319;
			18218: outdata = 32'd47318;
			18219: outdata = 32'd47317;
			18220: outdata = 32'd47316;
			18221: outdata = 32'd47315;
			18222: outdata = 32'd47314;
			18223: outdata = 32'd47313;
			18224: outdata = 32'd47312;
			18225: outdata = 32'd47311;
			18226: outdata = 32'd47310;
			18227: outdata = 32'd47309;
			18228: outdata = 32'd47308;
			18229: outdata = 32'd47307;
			18230: outdata = 32'd47306;
			18231: outdata = 32'd47305;
			18232: outdata = 32'd47304;
			18233: outdata = 32'd47303;
			18234: outdata = 32'd47302;
			18235: outdata = 32'd47301;
			18236: outdata = 32'd47300;
			18237: outdata = 32'd47299;
			18238: outdata = 32'd47298;
			18239: outdata = 32'd47297;
			18240: outdata = 32'd47296;
			18241: outdata = 32'd47295;
			18242: outdata = 32'd47294;
			18243: outdata = 32'd47293;
			18244: outdata = 32'd47292;
			18245: outdata = 32'd47291;
			18246: outdata = 32'd47290;
			18247: outdata = 32'd47289;
			18248: outdata = 32'd47288;
			18249: outdata = 32'd47287;
			18250: outdata = 32'd47286;
			18251: outdata = 32'd47285;
			18252: outdata = 32'd47284;
			18253: outdata = 32'd47283;
			18254: outdata = 32'd47282;
			18255: outdata = 32'd47281;
			18256: outdata = 32'd47280;
			18257: outdata = 32'd47279;
			18258: outdata = 32'd47278;
			18259: outdata = 32'd47277;
			18260: outdata = 32'd47276;
			18261: outdata = 32'd47275;
			18262: outdata = 32'd47274;
			18263: outdata = 32'd47273;
			18264: outdata = 32'd47272;
			18265: outdata = 32'd47271;
			18266: outdata = 32'd47270;
			18267: outdata = 32'd47269;
			18268: outdata = 32'd47268;
			18269: outdata = 32'd47267;
			18270: outdata = 32'd47266;
			18271: outdata = 32'd47265;
			18272: outdata = 32'd47264;
			18273: outdata = 32'd47263;
			18274: outdata = 32'd47262;
			18275: outdata = 32'd47261;
			18276: outdata = 32'd47260;
			18277: outdata = 32'd47259;
			18278: outdata = 32'd47258;
			18279: outdata = 32'd47257;
			18280: outdata = 32'd47256;
			18281: outdata = 32'd47255;
			18282: outdata = 32'd47254;
			18283: outdata = 32'd47253;
			18284: outdata = 32'd47252;
			18285: outdata = 32'd47251;
			18286: outdata = 32'd47250;
			18287: outdata = 32'd47249;
			18288: outdata = 32'd47248;
			18289: outdata = 32'd47247;
			18290: outdata = 32'd47246;
			18291: outdata = 32'd47245;
			18292: outdata = 32'd47244;
			18293: outdata = 32'd47243;
			18294: outdata = 32'd47242;
			18295: outdata = 32'd47241;
			18296: outdata = 32'd47240;
			18297: outdata = 32'd47239;
			18298: outdata = 32'd47238;
			18299: outdata = 32'd47237;
			18300: outdata = 32'd47236;
			18301: outdata = 32'd47235;
			18302: outdata = 32'd47234;
			18303: outdata = 32'd47233;
			18304: outdata = 32'd47232;
			18305: outdata = 32'd47231;
			18306: outdata = 32'd47230;
			18307: outdata = 32'd47229;
			18308: outdata = 32'd47228;
			18309: outdata = 32'd47227;
			18310: outdata = 32'd47226;
			18311: outdata = 32'd47225;
			18312: outdata = 32'd47224;
			18313: outdata = 32'd47223;
			18314: outdata = 32'd47222;
			18315: outdata = 32'd47221;
			18316: outdata = 32'd47220;
			18317: outdata = 32'd47219;
			18318: outdata = 32'd47218;
			18319: outdata = 32'd47217;
			18320: outdata = 32'd47216;
			18321: outdata = 32'd47215;
			18322: outdata = 32'd47214;
			18323: outdata = 32'd47213;
			18324: outdata = 32'd47212;
			18325: outdata = 32'd47211;
			18326: outdata = 32'd47210;
			18327: outdata = 32'd47209;
			18328: outdata = 32'd47208;
			18329: outdata = 32'd47207;
			18330: outdata = 32'd47206;
			18331: outdata = 32'd47205;
			18332: outdata = 32'd47204;
			18333: outdata = 32'd47203;
			18334: outdata = 32'd47202;
			18335: outdata = 32'd47201;
			18336: outdata = 32'd47200;
			18337: outdata = 32'd47199;
			18338: outdata = 32'd47198;
			18339: outdata = 32'd47197;
			18340: outdata = 32'd47196;
			18341: outdata = 32'd47195;
			18342: outdata = 32'd47194;
			18343: outdata = 32'd47193;
			18344: outdata = 32'd47192;
			18345: outdata = 32'd47191;
			18346: outdata = 32'd47190;
			18347: outdata = 32'd47189;
			18348: outdata = 32'd47188;
			18349: outdata = 32'd47187;
			18350: outdata = 32'd47186;
			18351: outdata = 32'd47185;
			18352: outdata = 32'd47184;
			18353: outdata = 32'd47183;
			18354: outdata = 32'd47182;
			18355: outdata = 32'd47181;
			18356: outdata = 32'd47180;
			18357: outdata = 32'd47179;
			18358: outdata = 32'd47178;
			18359: outdata = 32'd47177;
			18360: outdata = 32'd47176;
			18361: outdata = 32'd47175;
			18362: outdata = 32'd47174;
			18363: outdata = 32'd47173;
			18364: outdata = 32'd47172;
			18365: outdata = 32'd47171;
			18366: outdata = 32'd47170;
			18367: outdata = 32'd47169;
			18368: outdata = 32'd47168;
			18369: outdata = 32'd47167;
			18370: outdata = 32'd47166;
			18371: outdata = 32'd47165;
			18372: outdata = 32'd47164;
			18373: outdata = 32'd47163;
			18374: outdata = 32'd47162;
			18375: outdata = 32'd47161;
			18376: outdata = 32'd47160;
			18377: outdata = 32'd47159;
			18378: outdata = 32'd47158;
			18379: outdata = 32'd47157;
			18380: outdata = 32'd47156;
			18381: outdata = 32'd47155;
			18382: outdata = 32'd47154;
			18383: outdata = 32'd47153;
			18384: outdata = 32'd47152;
			18385: outdata = 32'd47151;
			18386: outdata = 32'd47150;
			18387: outdata = 32'd47149;
			18388: outdata = 32'd47148;
			18389: outdata = 32'd47147;
			18390: outdata = 32'd47146;
			18391: outdata = 32'd47145;
			18392: outdata = 32'd47144;
			18393: outdata = 32'd47143;
			18394: outdata = 32'd47142;
			18395: outdata = 32'd47141;
			18396: outdata = 32'd47140;
			18397: outdata = 32'd47139;
			18398: outdata = 32'd47138;
			18399: outdata = 32'd47137;
			18400: outdata = 32'd47136;
			18401: outdata = 32'd47135;
			18402: outdata = 32'd47134;
			18403: outdata = 32'd47133;
			18404: outdata = 32'd47132;
			18405: outdata = 32'd47131;
			18406: outdata = 32'd47130;
			18407: outdata = 32'd47129;
			18408: outdata = 32'd47128;
			18409: outdata = 32'd47127;
			18410: outdata = 32'd47126;
			18411: outdata = 32'd47125;
			18412: outdata = 32'd47124;
			18413: outdata = 32'd47123;
			18414: outdata = 32'd47122;
			18415: outdata = 32'd47121;
			18416: outdata = 32'd47120;
			18417: outdata = 32'd47119;
			18418: outdata = 32'd47118;
			18419: outdata = 32'd47117;
			18420: outdata = 32'd47116;
			18421: outdata = 32'd47115;
			18422: outdata = 32'd47114;
			18423: outdata = 32'd47113;
			18424: outdata = 32'd47112;
			18425: outdata = 32'd47111;
			18426: outdata = 32'd47110;
			18427: outdata = 32'd47109;
			18428: outdata = 32'd47108;
			18429: outdata = 32'd47107;
			18430: outdata = 32'd47106;
			18431: outdata = 32'd47105;
			18432: outdata = 32'd47104;
			18433: outdata = 32'd47103;
			18434: outdata = 32'd47102;
			18435: outdata = 32'd47101;
			18436: outdata = 32'd47100;
			18437: outdata = 32'd47099;
			18438: outdata = 32'd47098;
			18439: outdata = 32'd47097;
			18440: outdata = 32'd47096;
			18441: outdata = 32'd47095;
			18442: outdata = 32'd47094;
			18443: outdata = 32'd47093;
			18444: outdata = 32'd47092;
			18445: outdata = 32'd47091;
			18446: outdata = 32'd47090;
			18447: outdata = 32'd47089;
			18448: outdata = 32'd47088;
			18449: outdata = 32'd47087;
			18450: outdata = 32'd47086;
			18451: outdata = 32'd47085;
			18452: outdata = 32'd47084;
			18453: outdata = 32'd47083;
			18454: outdata = 32'd47082;
			18455: outdata = 32'd47081;
			18456: outdata = 32'd47080;
			18457: outdata = 32'd47079;
			18458: outdata = 32'd47078;
			18459: outdata = 32'd47077;
			18460: outdata = 32'd47076;
			18461: outdata = 32'd47075;
			18462: outdata = 32'd47074;
			18463: outdata = 32'd47073;
			18464: outdata = 32'd47072;
			18465: outdata = 32'd47071;
			18466: outdata = 32'd47070;
			18467: outdata = 32'd47069;
			18468: outdata = 32'd47068;
			18469: outdata = 32'd47067;
			18470: outdata = 32'd47066;
			18471: outdata = 32'd47065;
			18472: outdata = 32'd47064;
			18473: outdata = 32'd47063;
			18474: outdata = 32'd47062;
			18475: outdata = 32'd47061;
			18476: outdata = 32'd47060;
			18477: outdata = 32'd47059;
			18478: outdata = 32'd47058;
			18479: outdata = 32'd47057;
			18480: outdata = 32'd47056;
			18481: outdata = 32'd47055;
			18482: outdata = 32'd47054;
			18483: outdata = 32'd47053;
			18484: outdata = 32'd47052;
			18485: outdata = 32'd47051;
			18486: outdata = 32'd47050;
			18487: outdata = 32'd47049;
			18488: outdata = 32'd47048;
			18489: outdata = 32'd47047;
			18490: outdata = 32'd47046;
			18491: outdata = 32'd47045;
			18492: outdata = 32'd47044;
			18493: outdata = 32'd47043;
			18494: outdata = 32'd47042;
			18495: outdata = 32'd47041;
			18496: outdata = 32'd47040;
			18497: outdata = 32'd47039;
			18498: outdata = 32'd47038;
			18499: outdata = 32'd47037;
			18500: outdata = 32'd47036;
			18501: outdata = 32'd47035;
			18502: outdata = 32'd47034;
			18503: outdata = 32'd47033;
			18504: outdata = 32'd47032;
			18505: outdata = 32'd47031;
			18506: outdata = 32'd47030;
			18507: outdata = 32'd47029;
			18508: outdata = 32'd47028;
			18509: outdata = 32'd47027;
			18510: outdata = 32'd47026;
			18511: outdata = 32'd47025;
			18512: outdata = 32'd47024;
			18513: outdata = 32'd47023;
			18514: outdata = 32'd47022;
			18515: outdata = 32'd47021;
			18516: outdata = 32'd47020;
			18517: outdata = 32'd47019;
			18518: outdata = 32'd47018;
			18519: outdata = 32'd47017;
			18520: outdata = 32'd47016;
			18521: outdata = 32'd47015;
			18522: outdata = 32'd47014;
			18523: outdata = 32'd47013;
			18524: outdata = 32'd47012;
			18525: outdata = 32'd47011;
			18526: outdata = 32'd47010;
			18527: outdata = 32'd47009;
			18528: outdata = 32'd47008;
			18529: outdata = 32'd47007;
			18530: outdata = 32'd47006;
			18531: outdata = 32'd47005;
			18532: outdata = 32'd47004;
			18533: outdata = 32'd47003;
			18534: outdata = 32'd47002;
			18535: outdata = 32'd47001;
			18536: outdata = 32'd47000;
			18537: outdata = 32'd46999;
			18538: outdata = 32'd46998;
			18539: outdata = 32'd46997;
			18540: outdata = 32'd46996;
			18541: outdata = 32'd46995;
			18542: outdata = 32'd46994;
			18543: outdata = 32'd46993;
			18544: outdata = 32'd46992;
			18545: outdata = 32'd46991;
			18546: outdata = 32'd46990;
			18547: outdata = 32'd46989;
			18548: outdata = 32'd46988;
			18549: outdata = 32'd46987;
			18550: outdata = 32'd46986;
			18551: outdata = 32'd46985;
			18552: outdata = 32'd46984;
			18553: outdata = 32'd46983;
			18554: outdata = 32'd46982;
			18555: outdata = 32'd46981;
			18556: outdata = 32'd46980;
			18557: outdata = 32'd46979;
			18558: outdata = 32'd46978;
			18559: outdata = 32'd46977;
			18560: outdata = 32'd46976;
			18561: outdata = 32'd46975;
			18562: outdata = 32'd46974;
			18563: outdata = 32'd46973;
			18564: outdata = 32'd46972;
			18565: outdata = 32'd46971;
			18566: outdata = 32'd46970;
			18567: outdata = 32'd46969;
			18568: outdata = 32'd46968;
			18569: outdata = 32'd46967;
			18570: outdata = 32'd46966;
			18571: outdata = 32'd46965;
			18572: outdata = 32'd46964;
			18573: outdata = 32'd46963;
			18574: outdata = 32'd46962;
			18575: outdata = 32'd46961;
			18576: outdata = 32'd46960;
			18577: outdata = 32'd46959;
			18578: outdata = 32'd46958;
			18579: outdata = 32'd46957;
			18580: outdata = 32'd46956;
			18581: outdata = 32'd46955;
			18582: outdata = 32'd46954;
			18583: outdata = 32'd46953;
			18584: outdata = 32'd46952;
			18585: outdata = 32'd46951;
			18586: outdata = 32'd46950;
			18587: outdata = 32'd46949;
			18588: outdata = 32'd46948;
			18589: outdata = 32'd46947;
			18590: outdata = 32'd46946;
			18591: outdata = 32'd46945;
			18592: outdata = 32'd46944;
			18593: outdata = 32'd46943;
			18594: outdata = 32'd46942;
			18595: outdata = 32'd46941;
			18596: outdata = 32'd46940;
			18597: outdata = 32'd46939;
			18598: outdata = 32'd46938;
			18599: outdata = 32'd46937;
			18600: outdata = 32'd46936;
			18601: outdata = 32'd46935;
			18602: outdata = 32'd46934;
			18603: outdata = 32'd46933;
			18604: outdata = 32'd46932;
			18605: outdata = 32'd46931;
			18606: outdata = 32'd46930;
			18607: outdata = 32'd46929;
			18608: outdata = 32'd46928;
			18609: outdata = 32'd46927;
			18610: outdata = 32'd46926;
			18611: outdata = 32'd46925;
			18612: outdata = 32'd46924;
			18613: outdata = 32'd46923;
			18614: outdata = 32'd46922;
			18615: outdata = 32'd46921;
			18616: outdata = 32'd46920;
			18617: outdata = 32'd46919;
			18618: outdata = 32'd46918;
			18619: outdata = 32'd46917;
			18620: outdata = 32'd46916;
			18621: outdata = 32'd46915;
			18622: outdata = 32'd46914;
			18623: outdata = 32'd46913;
			18624: outdata = 32'd46912;
			18625: outdata = 32'd46911;
			18626: outdata = 32'd46910;
			18627: outdata = 32'd46909;
			18628: outdata = 32'd46908;
			18629: outdata = 32'd46907;
			18630: outdata = 32'd46906;
			18631: outdata = 32'd46905;
			18632: outdata = 32'd46904;
			18633: outdata = 32'd46903;
			18634: outdata = 32'd46902;
			18635: outdata = 32'd46901;
			18636: outdata = 32'd46900;
			18637: outdata = 32'd46899;
			18638: outdata = 32'd46898;
			18639: outdata = 32'd46897;
			18640: outdata = 32'd46896;
			18641: outdata = 32'd46895;
			18642: outdata = 32'd46894;
			18643: outdata = 32'd46893;
			18644: outdata = 32'd46892;
			18645: outdata = 32'd46891;
			18646: outdata = 32'd46890;
			18647: outdata = 32'd46889;
			18648: outdata = 32'd46888;
			18649: outdata = 32'd46887;
			18650: outdata = 32'd46886;
			18651: outdata = 32'd46885;
			18652: outdata = 32'd46884;
			18653: outdata = 32'd46883;
			18654: outdata = 32'd46882;
			18655: outdata = 32'd46881;
			18656: outdata = 32'd46880;
			18657: outdata = 32'd46879;
			18658: outdata = 32'd46878;
			18659: outdata = 32'd46877;
			18660: outdata = 32'd46876;
			18661: outdata = 32'd46875;
			18662: outdata = 32'd46874;
			18663: outdata = 32'd46873;
			18664: outdata = 32'd46872;
			18665: outdata = 32'd46871;
			18666: outdata = 32'd46870;
			18667: outdata = 32'd46869;
			18668: outdata = 32'd46868;
			18669: outdata = 32'd46867;
			18670: outdata = 32'd46866;
			18671: outdata = 32'd46865;
			18672: outdata = 32'd46864;
			18673: outdata = 32'd46863;
			18674: outdata = 32'd46862;
			18675: outdata = 32'd46861;
			18676: outdata = 32'd46860;
			18677: outdata = 32'd46859;
			18678: outdata = 32'd46858;
			18679: outdata = 32'd46857;
			18680: outdata = 32'd46856;
			18681: outdata = 32'd46855;
			18682: outdata = 32'd46854;
			18683: outdata = 32'd46853;
			18684: outdata = 32'd46852;
			18685: outdata = 32'd46851;
			18686: outdata = 32'd46850;
			18687: outdata = 32'd46849;
			18688: outdata = 32'd46848;
			18689: outdata = 32'd46847;
			18690: outdata = 32'd46846;
			18691: outdata = 32'd46845;
			18692: outdata = 32'd46844;
			18693: outdata = 32'd46843;
			18694: outdata = 32'd46842;
			18695: outdata = 32'd46841;
			18696: outdata = 32'd46840;
			18697: outdata = 32'd46839;
			18698: outdata = 32'd46838;
			18699: outdata = 32'd46837;
			18700: outdata = 32'd46836;
			18701: outdata = 32'd46835;
			18702: outdata = 32'd46834;
			18703: outdata = 32'd46833;
			18704: outdata = 32'd46832;
			18705: outdata = 32'd46831;
			18706: outdata = 32'd46830;
			18707: outdata = 32'd46829;
			18708: outdata = 32'd46828;
			18709: outdata = 32'd46827;
			18710: outdata = 32'd46826;
			18711: outdata = 32'd46825;
			18712: outdata = 32'd46824;
			18713: outdata = 32'd46823;
			18714: outdata = 32'd46822;
			18715: outdata = 32'd46821;
			18716: outdata = 32'd46820;
			18717: outdata = 32'd46819;
			18718: outdata = 32'd46818;
			18719: outdata = 32'd46817;
			18720: outdata = 32'd46816;
			18721: outdata = 32'd46815;
			18722: outdata = 32'd46814;
			18723: outdata = 32'd46813;
			18724: outdata = 32'd46812;
			18725: outdata = 32'd46811;
			18726: outdata = 32'd46810;
			18727: outdata = 32'd46809;
			18728: outdata = 32'd46808;
			18729: outdata = 32'd46807;
			18730: outdata = 32'd46806;
			18731: outdata = 32'd46805;
			18732: outdata = 32'd46804;
			18733: outdata = 32'd46803;
			18734: outdata = 32'd46802;
			18735: outdata = 32'd46801;
			18736: outdata = 32'd46800;
			18737: outdata = 32'd46799;
			18738: outdata = 32'd46798;
			18739: outdata = 32'd46797;
			18740: outdata = 32'd46796;
			18741: outdata = 32'd46795;
			18742: outdata = 32'd46794;
			18743: outdata = 32'd46793;
			18744: outdata = 32'd46792;
			18745: outdata = 32'd46791;
			18746: outdata = 32'd46790;
			18747: outdata = 32'd46789;
			18748: outdata = 32'd46788;
			18749: outdata = 32'd46787;
			18750: outdata = 32'd46786;
			18751: outdata = 32'd46785;
			18752: outdata = 32'd46784;
			18753: outdata = 32'd46783;
			18754: outdata = 32'd46782;
			18755: outdata = 32'd46781;
			18756: outdata = 32'd46780;
			18757: outdata = 32'd46779;
			18758: outdata = 32'd46778;
			18759: outdata = 32'd46777;
			18760: outdata = 32'd46776;
			18761: outdata = 32'd46775;
			18762: outdata = 32'd46774;
			18763: outdata = 32'd46773;
			18764: outdata = 32'd46772;
			18765: outdata = 32'd46771;
			18766: outdata = 32'd46770;
			18767: outdata = 32'd46769;
			18768: outdata = 32'd46768;
			18769: outdata = 32'd46767;
			18770: outdata = 32'd46766;
			18771: outdata = 32'd46765;
			18772: outdata = 32'd46764;
			18773: outdata = 32'd46763;
			18774: outdata = 32'd46762;
			18775: outdata = 32'd46761;
			18776: outdata = 32'd46760;
			18777: outdata = 32'd46759;
			18778: outdata = 32'd46758;
			18779: outdata = 32'd46757;
			18780: outdata = 32'd46756;
			18781: outdata = 32'd46755;
			18782: outdata = 32'd46754;
			18783: outdata = 32'd46753;
			18784: outdata = 32'd46752;
			18785: outdata = 32'd46751;
			18786: outdata = 32'd46750;
			18787: outdata = 32'd46749;
			18788: outdata = 32'd46748;
			18789: outdata = 32'd46747;
			18790: outdata = 32'd46746;
			18791: outdata = 32'd46745;
			18792: outdata = 32'd46744;
			18793: outdata = 32'd46743;
			18794: outdata = 32'd46742;
			18795: outdata = 32'd46741;
			18796: outdata = 32'd46740;
			18797: outdata = 32'd46739;
			18798: outdata = 32'd46738;
			18799: outdata = 32'd46737;
			18800: outdata = 32'd46736;
			18801: outdata = 32'd46735;
			18802: outdata = 32'd46734;
			18803: outdata = 32'd46733;
			18804: outdata = 32'd46732;
			18805: outdata = 32'd46731;
			18806: outdata = 32'd46730;
			18807: outdata = 32'd46729;
			18808: outdata = 32'd46728;
			18809: outdata = 32'd46727;
			18810: outdata = 32'd46726;
			18811: outdata = 32'd46725;
			18812: outdata = 32'd46724;
			18813: outdata = 32'd46723;
			18814: outdata = 32'd46722;
			18815: outdata = 32'd46721;
			18816: outdata = 32'd46720;
			18817: outdata = 32'd46719;
			18818: outdata = 32'd46718;
			18819: outdata = 32'd46717;
			18820: outdata = 32'd46716;
			18821: outdata = 32'd46715;
			18822: outdata = 32'd46714;
			18823: outdata = 32'd46713;
			18824: outdata = 32'd46712;
			18825: outdata = 32'd46711;
			18826: outdata = 32'd46710;
			18827: outdata = 32'd46709;
			18828: outdata = 32'd46708;
			18829: outdata = 32'd46707;
			18830: outdata = 32'd46706;
			18831: outdata = 32'd46705;
			18832: outdata = 32'd46704;
			18833: outdata = 32'd46703;
			18834: outdata = 32'd46702;
			18835: outdata = 32'd46701;
			18836: outdata = 32'd46700;
			18837: outdata = 32'd46699;
			18838: outdata = 32'd46698;
			18839: outdata = 32'd46697;
			18840: outdata = 32'd46696;
			18841: outdata = 32'd46695;
			18842: outdata = 32'd46694;
			18843: outdata = 32'd46693;
			18844: outdata = 32'd46692;
			18845: outdata = 32'd46691;
			18846: outdata = 32'd46690;
			18847: outdata = 32'd46689;
			18848: outdata = 32'd46688;
			18849: outdata = 32'd46687;
			18850: outdata = 32'd46686;
			18851: outdata = 32'd46685;
			18852: outdata = 32'd46684;
			18853: outdata = 32'd46683;
			18854: outdata = 32'd46682;
			18855: outdata = 32'd46681;
			18856: outdata = 32'd46680;
			18857: outdata = 32'd46679;
			18858: outdata = 32'd46678;
			18859: outdata = 32'd46677;
			18860: outdata = 32'd46676;
			18861: outdata = 32'd46675;
			18862: outdata = 32'd46674;
			18863: outdata = 32'd46673;
			18864: outdata = 32'd46672;
			18865: outdata = 32'd46671;
			18866: outdata = 32'd46670;
			18867: outdata = 32'd46669;
			18868: outdata = 32'd46668;
			18869: outdata = 32'd46667;
			18870: outdata = 32'd46666;
			18871: outdata = 32'd46665;
			18872: outdata = 32'd46664;
			18873: outdata = 32'd46663;
			18874: outdata = 32'd46662;
			18875: outdata = 32'd46661;
			18876: outdata = 32'd46660;
			18877: outdata = 32'd46659;
			18878: outdata = 32'd46658;
			18879: outdata = 32'd46657;
			18880: outdata = 32'd46656;
			18881: outdata = 32'd46655;
			18882: outdata = 32'd46654;
			18883: outdata = 32'd46653;
			18884: outdata = 32'd46652;
			18885: outdata = 32'd46651;
			18886: outdata = 32'd46650;
			18887: outdata = 32'd46649;
			18888: outdata = 32'd46648;
			18889: outdata = 32'd46647;
			18890: outdata = 32'd46646;
			18891: outdata = 32'd46645;
			18892: outdata = 32'd46644;
			18893: outdata = 32'd46643;
			18894: outdata = 32'd46642;
			18895: outdata = 32'd46641;
			18896: outdata = 32'd46640;
			18897: outdata = 32'd46639;
			18898: outdata = 32'd46638;
			18899: outdata = 32'd46637;
			18900: outdata = 32'd46636;
			18901: outdata = 32'd46635;
			18902: outdata = 32'd46634;
			18903: outdata = 32'd46633;
			18904: outdata = 32'd46632;
			18905: outdata = 32'd46631;
			18906: outdata = 32'd46630;
			18907: outdata = 32'd46629;
			18908: outdata = 32'd46628;
			18909: outdata = 32'd46627;
			18910: outdata = 32'd46626;
			18911: outdata = 32'd46625;
			18912: outdata = 32'd46624;
			18913: outdata = 32'd46623;
			18914: outdata = 32'd46622;
			18915: outdata = 32'd46621;
			18916: outdata = 32'd46620;
			18917: outdata = 32'd46619;
			18918: outdata = 32'd46618;
			18919: outdata = 32'd46617;
			18920: outdata = 32'd46616;
			18921: outdata = 32'd46615;
			18922: outdata = 32'd46614;
			18923: outdata = 32'd46613;
			18924: outdata = 32'd46612;
			18925: outdata = 32'd46611;
			18926: outdata = 32'd46610;
			18927: outdata = 32'd46609;
			18928: outdata = 32'd46608;
			18929: outdata = 32'd46607;
			18930: outdata = 32'd46606;
			18931: outdata = 32'd46605;
			18932: outdata = 32'd46604;
			18933: outdata = 32'd46603;
			18934: outdata = 32'd46602;
			18935: outdata = 32'd46601;
			18936: outdata = 32'd46600;
			18937: outdata = 32'd46599;
			18938: outdata = 32'd46598;
			18939: outdata = 32'd46597;
			18940: outdata = 32'd46596;
			18941: outdata = 32'd46595;
			18942: outdata = 32'd46594;
			18943: outdata = 32'd46593;
			18944: outdata = 32'd46592;
			18945: outdata = 32'd46591;
			18946: outdata = 32'd46590;
			18947: outdata = 32'd46589;
			18948: outdata = 32'd46588;
			18949: outdata = 32'd46587;
			18950: outdata = 32'd46586;
			18951: outdata = 32'd46585;
			18952: outdata = 32'd46584;
			18953: outdata = 32'd46583;
			18954: outdata = 32'd46582;
			18955: outdata = 32'd46581;
			18956: outdata = 32'd46580;
			18957: outdata = 32'd46579;
			18958: outdata = 32'd46578;
			18959: outdata = 32'd46577;
			18960: outdata = 32'd46576;
			18961: outdata = 32'd46575;
			18962: outdata = 32'd46574;
			18963: outdata = 32'd46573;
			18964: outdata = 32'd46572;
			18965: outdata = 32'd46571;
			18966: outdata = 32'd46570;
			18967: outdata = 32'd46569;
			18968: outdata = 32'd46568;
			18969: outdata = 32'd46567;
			18970: outdata = 32'd46566;
			18971: outdata = 32'd46565;
			18972: outdata = 32'd46564;
			18973: outdata = 32'd46563;
			18974: outdata = 32'd46562;
			18975: outdata = 32'd46561;
			18976: outdata = 32'd46560;
			18977: outdata = 32'd46559;
			18978: outdata = 32'd46558;
			18979: outdata = 32'd46557;
			18980: outdata = 32'd46556;
			18981: outdata = 32'd46555;
			18982: outdata = 32'd46554;
			18983: outdata = 32'd46553;
			18984: outdata = 32'd46552;
			18985: outdata = 32'd46551;
			18986: outdata = 32'd46550;
			18987: outdata = 32'd46549;
			18988: outdata = 32'd46548;
			18989: outdata = 32'd46547;
			18990: outdata = 32'd46546;
			18991: outdata = 32'd46545;
			18992: outdata = 32'd46544;
			18993: outdata = 32'd46543;
			18994: outdata = 32'd46542;
			18995: outdata = 32'd46541;
			18996: outdata = 32'd46540;
			18997: outdata = 32'd46539;
			18998: outdata = 32'd46538;
			18999: outdata = 32'd46537;
			19000: outdata = 32'd46536;
			19001: outdata = 32'd46535;
			19002: outdata = 32'd46534;
			19003: outdata = 32'd46533;
			19004: outdata = 32'd46532;
			19005: outdata = 32'd46531;
			19006: outdata = 32'd46530;
			19007: outdata = 32'd46529;
			19008: outdata = 32'd46528;
			19009: outdata = 32'd46527;
			19010: outdata = 32'd46526;
			19011: outdata = 32'd46525;
			19012: outdata = 32'd46524;
			19013: outdata = 32'd46523;
			19014: outdata = 32'd46522;
			19015: outdata = 32'd46521;
			19016: outdata = 32'd46520;
			19017: outdata = 32'd46519;
			19018: outdata = 32'd46518;
			19019: outdata = 32'd46517;
			19020: outdata = 32'd46516;
			19021: outdata = 32'd46515;
			19022: outdata = 32'd46514;
			19023: outdata = 32'd46513;
			19024: outdata = 32'd46512;
			19025: outdata = 32'd46511;
			19026: outdata = 32'd46510;
			19027: outdata = 32'd46509;
			19028: outdata = 32'd46508;
			19029: outdata = 32'd46507;
			19030: outdata = 32'd46506;
			19031: outdata = 32'd46505;
			19032: outdata = 32'd46504;
			19033: outdata = 32'd46503;
			19034: outdata = 32'd46502;
			19035: outdata = 32'd46501;
			19036: outdata = 32'd46500;
			19037: outdata = 32'd46499;
			19038: outdata = 32'd46498;
			19039: outdata = 32'd46497;
			19040: outdata = 32'd46496;
			19041: outdata = 32'd46495;
			19042: outdata = 32'd46494;
			19043: outdata = 32'd46493;
			19044: outdata = 32'd46492;
			19045: outdata = 32'd46491;
			19046: outdata = 32'd46490;
			19047: outdata = 32'd46489;
			19048: outdata = 32'd46488;
			19049: outdata = 32'd46487;
			19050: outdata = 32'd46486;
			19051: outdata = 32'd46485;
			19052: outdata = 32'd46484;
			19053: outdata = 32'd46483;
			19054: outdata = 32'd46482;
			19055: outdata = 32'd46481;
			19056: outdata = 32'd46480;
			19057: outdata = 32'd46479;
			19058: outdata = 32'd46478;
			19059: outdata = 32'd46477;
			19060: outdata = 32'd46476;
			19061: outdata = 32'd46475;
			19062: outdata = 32'd46474;
			19063: outdata = 32'd46473;
			19064: outdata = 32'd46472;
			19065: outdata = 32'd46471;
			19066: outdata = 32'd46470;
			19067: outdata = 32'd46469;
			19068: outdata = 32'd46468;
			19069: outdata = 32'd46467;
			19070: outdata = 32'd46466;
			19071: outdata = 32'd46465;
			19072: outdata = 32'd46464;
			19073: outdata = 32'd46463;
			19074: outdata = 32'd46462;
			19075: outdata = 32'd46461;
			19076: outdata = 32'd46460;
			19077: outdata = 32'd46459;
			19078: outdata = 32'd46458;
			19079: outdata = 32'd46457;
			19080: outdata = 32'd46456;
			19081: outdata = 32'd46455;
			19082: outdata = 32'd46454;
			19083: outdata = 32'd46453;
			19084: outdata = 32'd46452;
			19085: outdata = 32'd46451;
			19086: outdata = 32'd46450;
			19087: outdata = 32'd46449;
			19088: outdata = 32'd46448;
			19089: outdata = 32'd46447;
			19090: outdata = 32'd46446;
			19091: outdata = 32'd46445;
			19092: outdata = 32'd46444;
			19093: outdata = 32'd46443;
			19094: outdata = 32'd46442;
			19095: outdata = 32'd46441;
			19096: outdata = 32'd46440;
			19097: outdata = 32'd46439;
			19098: outdata = 32'd46438;
			19099: outdata = 32'd46437;
			19100: outdata = 32'd46436;
			19101: outdata = 32'd46435;
			19102: outdata = 32'd46434;
			19103: outdata = 32'd46433;
			19104: outdata = 32'd46432;
			19105: outdata = 32'd46431;
			19106: outdata = 32'd46430;
			19107: outdata = 32'd46429;
			19108: outdata = 32'd46428;
			19109: outdata = 32'd46427;
			19110: outdata = 32'd46426;
			19111: outdata = 32'd46425;
			19112: outdata = 32'd46424;
			19113: outdata = 32'd46423;
			19114: outdata = 32'd46422;
			19115: outdata = 32'd46421;
			19116: outdata = 32'd46420;
			19117: outdata = 32'd46419;
			19118: outdata = 32'd46418;
			19119: outdata = 32'd46417;
			19120: outdata = 32'd46416;
			19121: outdata = 32'd46415;
			19122: outdata = 32'd46414;
			19123: outdata = 32'd46413;
			19124: outdata = 32'd46412;
			19125: outdata = 32'd46411;
			19126: outdata = 32'd46410;
			19127: outdata = 32'd46409;
			19128: outdata = 32'd46408;
			19129: outdata = 32'd46407;
			19130: outdata = 32'd46406;
			19131: outdata = 32'd46405;
			19132: outdata = 32'd46404;
			19133: outdata = 32'd46403;
			19134: outdata = 32'd46402;
			19135: outdata = 32'd46401;
			19136: outdata = 32'd46400;
			19137: outdata = 32'd46399;
			19138: outdata = 32'd46398;
			19139: outdata = 32'd46397;
			19140: outdata = 32'd46396;
			19141: outdata = 32'd46395;
			19142: outdata = 32'd46394;
			19143: outdata = 32'd46393;
			19144: outdata = 32'd46392;
			19145: outdata = 32'd46391;
			19146: outdata = 32'd46390;
			19147: outdata = 32'd46389;
			19148: outdata = 32'd46388;
			19149: outdata = 32'd46387;
			19150: outdata = 32'd46386;
			19151: outdata = 32'd46385;
			19152: outdata = 32'd46384;
			19153: outdata = 32'd46383;
			19154: outdata = 32'd46382;
			19155: outdata = 32'd46381;
			19156: outdata = 32'd46380;
			19157: outdata = 32'd46379;
			19158: outdata = 32'd46378;
			19159: outdata = 32'd46377;
			19160: outdata = 32'd46376;
			19161: outdata = 32'd46375;
			19162: outdata = 32'd46374;
			19163: outdata = 32'd46373;
			19164: outdata = 32'd46372;
			19165: outdata = 32'd46371;
			19166: outdata = 32'd46370;
			19167: outdata = 32'd46369;
			19168: outdata = 32'd46368;
			19169: outdata = 32'd46367;
			19170: outdata = 32'd46366;
			19171: outdata = 32'd46365;
			19172: outdata = 32'd46364;
			19173: outdata = 32'd46363;
			19174: outdata = 32'd46362;
			19175: outdata = 32'd46361;
			19176: outdata = 32'd46360;
			19177: outdata = 32'd46359;
			19178: outdata = 32'd46358;
			19179: outdata = 32'd46357;
			19180: outdata = 32'd46356;
			19181: outdata = 32'd46355;
			19182: outdata = 32'd46354;
			19183: outdata = 32'd46353;
			19184: outdata = 32'd46352;
			19185: outdata = 32'd46351;
			19186: outdata = 32'd46350;
			19187: outdata = 32'd46349;
			19188: outdata = 32'd46348;
			19189: outdata = 32'd46347;
			19190: outdata = 32'd46346;
			19191: outdata = 32'd46345;
			19192: outdata = 32'd46344;
			19193: outdata = 32'd46343;
			19194: outdata = 32'd46342;
			19195: outdata = 32'd46341;
			19196: outdata = 32'd46340;
			19197: outdata = 32'd46339;
			19198: outdata = 32'd46338;
			19199: outdata = 32'd46337;
			19200: outdata = 32'd46336;
			19201: outdata = 32'd46335;
			19202: outdata = 32'd46334;
			19203: outdata = 32'd46333;
			19204: outdata = 32'd46332;
			19205: outdata = 32'd46331;
			19206: outdata = 32'd46330;
			19207: outdata = 32'd46329;
			19208: outdata = 32'd46328;
			19209: outdata = 32'd46327;
			19210: outdata = 32'd46326;
			19211: outdata = 32'd46325;
			19212: outdata = 32'd46324;
			19213: outdata = 32'd46323;
			19214: outdata = 32'd46322;
			19215: outdata = 32'd46321;
			19216: outdata = 32'd46320;
			19217: outdata = 32'd46319;
			19218: outdata = 32'd46318;
			19219: outdata = 32'd46317;
			19220: outdata = 32'd46316;
			19221: outdata = 32'd46315;
			19222: outdata = 32'd46314;
			19223: outdata = 32'd46313;
			19224: outdata = 32'd46312;
			19225: outdata = 32'd46311;
			19226: outdata = 32'd46310;
			19227: outdata = 32'd46309;
			19228: outdata = 32'd46308;
			19229: outdata = 32'd46307;
			19230: outdata = 32'd46306;
			19231: outdata = 32'd46305;
			19232: outdata = 32'd46304;
			19233: outdata = 32'd46303;
			19234: outdata = 32'd46302;
			19235: outdata = 32'd46301;
			19236: outdata = 32'd46300;
			19237: outdata = 32'd46299;
			19238: outdata = 32'd46298;
			19239: outdata = 32'd46297;
			19240: outdata = 32'd46296;
			19241: outdata = 32'd46295;
			19242: outdata = 32'd46294;
			19243: outdata = 32'd46293;
			19244: outdata = 32'd46292;
			19245: outdata = 32'd46291;
			19246: outdata = 32'd46290;
			19247: outdata = 32'd46289;
			19248: outdata = 32'd46288;
			19249: outdata = 32'd46287;
			19250: outdata = 32'd46286;
			19251: outdata = 32'd46285;
			19252: outdata = 32'd46284;
			19253: outdata = 32'd46283;
			19254: outdata = 32'd46282;
			19255: outdata = 32'd46281;
			19256: outdata = 32'd46280;
			19257: outdata = 32'd46279;
			19258: outdata = 32'd46278;
			19259: outdata = 32'd46277;
			19260: outdata = 32'd46276;
			19261: outdata = 32'd46275;
			19262: outdata = 32'd46274;
			19263: outdata = 32'd46273;
			19264: outdata = 32'd46272;
			19265: outdata = 32'd46271;
			19266: outdata = 32'd46270;
			19267: outdata = 32'd46269;
			19268: outdata = 32'd46268;
			19269: outdata = 32'd46267;
			19270: outdata = 32'd46266;
			19271: outdata = 32'd46265;
			19272: outdata = 32'd46264;
			19273: outdata = 32'd46263;
			19274: outdata = 32'd46262;
			19275: outdata = 32'd46261;
			19276: outdata = 32'd46260;
			19277: outdata = 32'd46259;
			19278: outdata = 32'd46258;
			19279: outdata = 32'd46257;
			19280: outdata = 32'd46256;
			19281: outdata = 32'd46255;
			19282: outdata = 32'd46254;
			19283: outdata = 32'd46253;
			19284: outdata = 32'd46252;
			19285: outdata = 32'd46251;
			19286: outdata = 32'd46250;
			19287: outdata = 32'd46249;
			19288: outdata = 32'd46248;
			19289: outdata = 32'd46247;
			19290: outdata = 32'd46246;
			19291: outdata = 32'd46245;
			19292: outdata = 32'd46244;
			19293: outdata = 32'd46243;
			19294: outdata = 32'd46242;
			19295: outdata = 32'd46241;
			19296: outdata = 32'd46240;
			19297: outdata = 32'd46239;
			19298: outdata = 32'd46238;
			19299: outdata = 32'd46237;
			19300: outdata = 32'd46236;
			19301: outdata = 32'd46235;
			19302: outdata = 32'd46234;
			19303: outdata = 32'd46233;
			19304: outdata = 32'd46232;
			19305: outdata = 32'd46231;
			19306: outdata = 32'd46230;
			19307: outdata = 32'd46229;
			19308: outdata = 32'd46228;
			19309: outdata = 32'd46227;
			19310: outdata = 32'd46226;
			19311: outdata = 32'd46225;
			19312: outdata = 32'd46224;
			19313: outdata = 32'd46223;
			19314: outdata = 32'd46222;
			19315: outdata = 32'd46221;
			19316: outdata = 32'd46220;
			19317: outdata = 32'd46219;
			19318: outdata = 32'd46218;
			19319: outdata = 32'd46217;
			19320: outdata = 32'd46216;
			19321: outdata = 32'd46215;
			19322: outdata = 32'd46214;
			19323: outdata = 32'd46213;
			19324: outdata = 32'd46212;
			19325: outdata = 32'd46211;
			19326: outdata = 32'd46210;
			19327: outdata = 32'd46209;
			19328: outdata = 32'd46208;
			19329: outdata = 32'd46207;
			19330: outdata = 32'd46206;
			19331: outdata = 32'd46205;
			19332: outdata = 32'd46204;
			19333: outdata = 32'd46203;
			19334: outdata = 32'd46202;
			19335: outdata = 32'd46201;
			19336: outdata = 32'd46200;
			19337: outdata = 32'd46199;
			19338: outdata = 32'd46198;
			19339: outdata = 32'd46197;
			19340: outdata = 32'd46196;
			19341: outdata = 32'd46195;
			19342: outdata = 32'd46194;
			19343: outdata = 32'd46193;
			19344: outdata = 32'd46192;
			19345: outdata = 32'd46191;
			19346: outdata = 32'd46190;
			19347: outdata = 32'd46189;
			19348: outdata = 32'd46188;
			19349: outdata = 32'd46187;
			19350: outdata = 32'd46186;
			19351: outdata = 32'd46185;
			19352: outdata = 32'd46184;
			19353: outdata = 32'd46183;
			19354: outdata = 32'd46182;
			19355: outdata = 32'd46181;
			19356: outdata = 32'd46180;
			19357: outdata = 32'd46179;
			19358: outdata = 32'd46178;
			19359: outdata = 32'd46177;
			19360: outdata = 32'd46176;
			19361: outdata = 32'd46175;
			19362: outdata = 32'd46174;
			19363: outdata = 32'd46173;
			19364: outdata = 32'd46172;
			19365: outdata = 32'd46171;
			19366: outdata = 32'd46170;
			19367: outdata = 32'd46169;
			19368: outdata = 32'd46168;
			19369: outdata = 32'd46167;
			19370: outdata = 32'd46166;
			19371: outdata = 32'd46165;
			19372: outdata = 32'd46164;
			19373: outdata = 32'd46163;
			19374: outdata = 32'd46162;
			19375: outdata = 32'd46161;
			19376: outdata = 32'd46160;
			19377: outdata = 32'd46159;
			19378: outdata = 32'd46158;
			19379: outdata = 32'd46157;
			19380: outdata = 32'd46156;
			19381: outdata = 32'd46155;
			19382: outdata = 32'd46154;
			19383: outdata = 32'd46153;
			19384: outdata = 32'd46152;
			19385: outdata = 32'd46151;
			19386: outdata = 32'd46150;
			19387: outdata = 32'd46149;
			19388: outdata = 32'd46148;
			19389: outdata = 32'd46147;
			19390: outdata = 32'd46146;
			19391: outdata = 32'd46145;
			19392: outdata = 32'd46144;
			19393: outdata = 32'd46143;
			19394: outdata = 32'd46142;
			19395: outdata = 32'd46141;
			19396: outdata = 32'd46140;
			19397: outdata = 32'd46139;
			19398: outdata = 32'd46138;
			19399: outdata = 32'd46137;
			19400: outdata = 32'd46136;
			19401: outdata = 32'd46135;
			19402: outdata = 32'd46134;
			19403: outdata = 32'd46133;
			19404: outdata = 32'd46132;
			19405: outdata = 32'd46131;
			19406: outdata = 32'd46130;
			19407: outdata = 32'd46129;
			19408: outdata = 32'd46128;
			19409: outdata = 32'd46127;
			19410: outdata = 32'd46126;
			19411: outdata = 32'd46125;
			19412: outdata = 32'd46124;
			19413: outdata = 32'd46123;
			19414: outdata = 32'd46122;
			19415: outdata = 32'd46121;
			19416: outdata = 32'd46120;
			19417: outdata = 32'd46119;
			19418: outdata = 32'd46118;
			19419: outdata = 32'd46117;
			19420: outdata = 32'd46116;
			19421: outdata = 32'd46115;
			19422: outdata = 32'd46114;
			19423: outdata = 32'd46113;
			19424: outdata = 32'd46112;
			19425: outdata = 32'd46111;
			19426: outdata = 32'd46110;
			19427: outdata = 32'd46109;
			19428: outdata = 32'd46108;
			19429: outdata = 32'd46107;
			19430: outdata = 32'd46106;
			19431: outdata = 32'd46105;
			19432: outdata = 32'd46104;
			19433: outdata = 32'd46103;
			19434: outdata = 32'd46102;
			19435: outdata = 32'd46101;
			19436: outdata = 32'd46100;
			19437: outdata = 32'd46099;
			19438: outdata = 32'd46098;
			19439: outdata = 32'd46097;
			19440: outdata = 32'd46096;
			19441: outdata = 32'd46095;
			19442: outdata = 32'd46094;
			19443: outdata = 32'd46093;
			19444: outdata = 32'd46092;
			19445: outdata = 32'd46091;
			19446: outdata = 32'd46090;
			19447: outdata = 32'd46089;
			19448: outdata = 32'd46088;
			19449: outdata = 32'd46087;
			19450: outdata = 32'd46086;
			19451: outdata = 32'd46085;
			19452: outdata = 32'd46084;
			19453: outdata = 32'd46083;
			19454: outdata = 32'd46082;
			19455: outdata = 32'd46081;
			19456: outdata = 32'd46080;
			19457: outdata = 32'd46079;
			19458: outdata = 32'd46078;
			19459: outdata = 32'd46077;
			19460: outdata = 32'd46076;
			19461: outdata = 32'd46075;
			19462: outdata = 32'd46074;
			19463: outdata = 32'd46073;
			19464: outdata = 32'd46072;
			19465: outdata = 32'd46071;
			19466: outdata = 32'd46070;
			19467: outdata = 32'd46069;
			19468: outdata = 32'd46068;
			19469: outdata = 32'd46067;
			19470: outdata = 32'd46066;
			19471: outdata = 32'd46065;
			19472: outdata = 32'd46064;
			19473: outdata = 32'd46063;
			19474: outdata = 32'd46062;
			19475: outdata = 32'd46061;
			19476: outdata = 32'd46060;
			19477: outdata = 32'd46059;
			19478: outdata = 32'd46058;
			19479: outdata = 32'd46057;
			19480: outdata = 32'd46056;
			19481: outdata = 32'd46055;
			19482: outdata = 32'd46054;
			19483: outdata = 32'd46053;
			19484: outdata = 32'd46052;
			19485: outdata = 32'd46051;
			19486: outdata = 32'd46050;
			19487: outdata = 32'd46049;
			19488: outdata = 32'd46048;
			19489: outdata = 32'd46047;
			19490: outdata = 32'd46046;
			19491: outdata = 32'd46045;
			19492: outdata = 32'd46044;
			19493: outdata = 32'd46043;
			19494: outdata = 32'd46042;
			19495: outdata = 32'd46041;
			19496: outdata = 32'd46040;
			19497: outdata = 32'd46039;
			19498: outdata = 32'd46038;
			19499: outdata = 32'd46037;
			19500: outdata = 32'd46036;
			19501: outdata = 32'd46035;
			19502: outdata = 32'd46034;
			19503: outdata = 32'd46033;
			19504: outdata = 32'd46032;
			19505: outdata = 32'd46031;
			19506: outdata = 32'd46030;
			19507: outdata = 32'd46029;
			19508: outdata = 32'd46028;
			19509: outdata = 32'd46027;
			19510: outdata = 32'd46026;
			19511: outdata = 32'd46025;
			19512: outdata = 32'd46024;
			19513: outdata = 32'd46023;
			19514: outdata = 32'd46022;
			19515: outdata = 32'd46021;
			19516: outdata = 32'd46020;
			19517: outdata = 32'd46019;
			19518: outdata = 32'd46018;
			19519: outdata = 32'd46017;
			19520: outdata = 32'd46016;
			19521: outdata = 32'd46015;
			19522: outdata = 32'd46014;
			19523: outdata = 32'd46013;
			19524: outdata = 32'd46012;
			19525: outdata = 32'd46011;
			19526: outdata = 32'd46010;
			19527: outdata = 32'd46009;
			19528: outdata = 32'd46008;
			19529: outdata = 32'd46007;
			19530: outdata = 32'd46006;
			19531: outdata = 32'd46005;
			19532: outdata = 32'd46004;
			19533: outdata = 32'd46003;
			19534: outdata = 32'd46002;
			19535: outdata = 32'd46001;
			19536: outdata = 32'd46000;
			19537: outdata = 32'd45999;
			19538: outdata = 32'd45998;
			19539: outdata = 32'd45997;
			19540: outdata = 32'd45996;
			19541: outdata = 32'd45995;
			19542: outdata = 32'd45994;
			19543: outdata = 32'd45993;
			19544: outdata = 32'd45992;
			19545: outdata = 32'd45991;
			19546: outdata = 32'd45990;
			19547: outdata = 32'd45989;
			19548: outdata = 32'd45988;
			19549: outdata = 32'd45987;
			19550: outdata = 32'd45986;
			19551: outdata = 32'd45985;
			19552: outdata = 32'd45984;
			19553: outdata = 32'd45983;
			19554: outdata = 32'd45982;
			19555: outdata = 32'd45981;
			19556: outdata = 32'd45980;
			19557: outdata = 32'd45979;
			19558: outdata = 32'd45978;
			19559: outdata = 32'd45977;
			19560: outdata = 32'd45976;
			19561: outdata = 32'd45975;
			19562: outdata = 32'd45974;
			19563: outdata = 32'd45973;
			19564: outdata = 32'd45972;
			19565: outdata = 32'd45971;
			19566: outdata = 32'd45970;
			19567: outdata = 32'd45969;
			19568: outdata = 32'd45968;
			19569: outdata = 32'd45967;
			19570: outdata = 32'd45966;
			19571: outdata = 32'd45965;
			19572: outdata = 32'd45964;
			19573: outdata = 32'd45963;
			19574: outdata = 32'd45962;
			19575: outdata = 32'd45961;
			19576: outdata = 32'd45960;
			19577: outdata = 32'd45959;
			19578: outdata = 32'd45958;
			19579: outdata = 32'd45957;
			19580: outdata = 32'd45956;
			19581: outdata = 32'd45955;
			19582: outdata = 32'd45954;
			19583: outdata = 32'd45953;
			19584: outdata = 32'd45952;
			19585: outdata = 32'd45951;
			19586: outdata = 32'd45950;
			19587: outdata = 32'd45949;
			19588: outdata = 32'd45948;
			19589: outdata = 32'd45947;
			19590: outdata = 32'd45946;
			19591: outdata = 32'd45945;
			19592: outdata = 32'd45944;
			19593: outdata = 32'd45943;
			19594: outdata = 32'd45942;
			19595: outdata = 32'd45941;
			19596: outdata = 32'd45940;
			19597: outdata = 32'd45939;
			19598: outdata = 32'd45938;
			19599: outdata = 32'd45937;
			19600: outdata = 32'd45936;
			19601: outdata = 32'd45935;
			19602: outdata = 32'd45934;
			19603: outdata = 32'd45933;
			19604: outdata = 32'd45932;
			19605: outdata = 32'd45931;
			19606: outdata = 32'd45930;
			19607: outdata = 32'd45929;
			19608: outdata = 32'd45928;
			19609: outdata = 32'd45927;
			19610: outdata = 32'd45926;
			19611: outdata = 32'd45925;
			19612: outdata = 32'd45924;
			19613: outdata = 32'd45923;
			19614: outdata = 32'd45922;
			19615: outdata = 32'd45921;
			19616: outdata = 32'd45920;
			19617: outdata = 32'd45919;
			19618: outdata = 32'd45918;
			19619: outdata = 32'd45917;
			19620: outdata = 32'd45916;
			19621: outdata = 32'd45915;
			19622: outdata = 32'd45914;
			19623: outdata = 32'd45913;
			19624: outdata = 32'd45912;
			19625: outdata = 32'd45911;
			19626: outdata = 32'd45910;
			19627: outdata = 32'd45909;
			19628: outdata = 32'd45908;
			19629: outdata = 32'd45907;
			19630: outdata = 32'd45906;
			19631: outdata = 32'd45905;
			19632: outdata = 32'd45904;
			19633: outdata = 32'd45903;
			19634: outdata = 32'd45902;
			19635: outdata = 32'd45901;
			19636: outdata = 32'd45900;
			19637: outdata = 32'd45899;
			19638: outdata = 32'd45898;
			19639: outdata = 32'd45897;
			19640: outdata = 32'd45896;
			19641: outdata = 32'd45895;
			19642: outdata = 32'd45894;
			19643: outdata = 32'd45893;
			19644: outdata = 32'd45892;
			19645: outdata = 32'd45891;
			19646: outdata = 32'd45890;
			19647: outdata = 32'd45889;
			19648: outdata = 32'd45888;
			19649: outdata = 32'd45887;
			19650: outdata = 32'd45886;
			19651: outdata = 32'd45885;
			19652: outdata = 32'd45884;
			19653: outdata = 32'd45883;
			19654: outdata = 32'd45882;
			19655: outdata = 32'd45881;
			19656: outdata = 32'd45880;
			19657: outdata = 32'd45879;
			19658: outdata = 32'd45878;
			19659: outdata = 32'd45877;
			19660: outdata = 32'd45876;
			19661: outdata = 32'd45875;
			19662: outdata = 32'd45874;
			19663: outdata = 32'd45873;
			19664: outdata = 32'd45872;
			19665: outdata = 32'd45871;
			19666: outdata = 32'd45870;
			19667: outdata = 32'd45869;
			19668: outdata = 32'd45868;
			19669: outdata = 32'd45867;
			19670: outdata = 32'd45866;
			19671: outdata = 32'd45865;
			19672: outdata = 32'd45864;
			19673: outdata = 32'd45863;
			19674: outdata = 32'd45862;
			19675: outdata = 32'd45861;
			19676: outdata = 32'd45860;
			19677: outdata = 32'd45859;
			19678: outdata = 32'd45858;
			19679: outdata = 32'd45857;
			19680: outdata = 32'd45856;
			19681: outdata = 32'd45855;
			19682: outdata = 32'd45854;
			19683: outdata = 32'd45853;
			19684: outdata = 32'd45852;
			19685: outdata = 32'd45851;
			19686: outdata = 32'd45850;
			19687: outdata = 32'd45849;
			19688: outdata = 32'd45848;
			19689: outdata = 32'd45847;
			19690: outdata = 32'd45846;
			19691: outdata = 32'd45845;
			19692: outdata = 32'd45844;
			19693: outdata = 32'd45843;
			19694: outdata = 32'd45842;
			19695: outdata = 32'd45841;
			19696: outdata = 32'd45840;
			19697: outdata = 32'd45839;
			19698: outdata = 32'd45838;
			19699: outdata = 32'd45837;
			19700: outdata = 32'd45836;
			19701: outdata = 32'd45835;
			19702: outdata = 32'd45834;
			19703: outdata = 32'd45833;
			19704: outdata = 32'd45832;
			19705: outdata = 32'd45831;
			19706: outdata = 32'd45830;
			19707: outdata = 32'd45829;
			19708: outdata = 32'd45828;
			19709: outdata = 32'd45827;
			19710: outdata = 32'd45826;
			19711: outdata = 32'd45825;
			19712: outdata = 32'd45824;
			19713: outdata = 32'd45823;
			19714: outdata = 32'd45822;
			19715: outdata = 32'd45821;
			19716: outdata = 32'd45820;
			19717: outdata = 32'd45819;
			19718: outdata = 32'd45818;
			19719: outdata = 32'd45817;
			19720: outdata = 32'd45816;
			19721: outdata = 32'd45815;
			19722: outdata = 32'd45814;
			19723: outdata = 32'd45813;
			19724: outdata = 32'd45812;
			19725: outdata = 32'd45811;
			19726: outdata = 32'd45810;
			19727: outdata = 32'd45809;
			19728: outdata = 32'd45808;
			19729: outdata = 32'd45807;
			19730: outdata = 32'd45806;
			19731: outdata = 32'd45805;
			19732: outdata = 32'd45804;
			19733: outdata = 32'd45803;
			19734: outdata = 32'd45802;
			19735: outdata = 32'd45801;
			19736: outdata = 32'd45800;
			19737: outdata = 32'd45799;
			19738: outdata = 32'd45798;
			19739: outdata = 32'd45797;
			19740: outdata = 32'd45796;
			19741: outdata = 32'd45795;
			19742: outdata = 32'd45794;
			19743: outdata = 32'd45793;
			19744: outdata = 32'd45792;
			19745: outdata = 32'd45791;
			19746: outdata = 32'd45790;
			19747: outdata = 32'd45789;
			19748: outdata = 32'd45788;
			19749: outdata = 32'd45787;
			19750: outdata = 32'd45786;
			19751: outdata = 32'd45785;
			19752: outdata = 32'd45784;
			19753: outdata = 32'd45783;
			19754: outdata = 32'd45782;
			19755: outdata = 32'd45781;
			19756: outdata = 32'd45780;
			19757: outdata = 32'd45779;
			19758: outdata = 32'd45778;
			19759: outdata = 32'd45777;
			19760: outdata = 32'd45776;
			19761: outdata = 32'd45775;
			19762: outdata = 32'd45774;
			19763: outdata = 32'd45773;
			19764: outdata = 32'd45772;
			19765: outdata = 32'd45771;
			19766: outdata = 32'd45770;
			19767: outdata = 32'd45769;
			19768: outdata = 32'd45768;
			19769: outdata = 32'd45767;
			19770: outdata = 32'd45766;
			19771: outdata = 32'd45765;
			19772: outdata = 32'd45764;
			19773: outdata = 32'd45763;
			19774: outdata = 32'd45762;
			19775: outdata = 32'd45761;
			19776: outdata = 32'd45760;
			19777: outdata = 32'd45759;
			19778: outdata = 32'd45758;
			19779: outdata = 32'd45757;
			19780: outdata = 32'd45756;
			19781: outdata = 32'd45755;
			19782: outdata = 32'd45754;
			19783: outdata = 32'd45753;
			19784: outdata = 32'd45752;
			19785: outdata = 32'd45751;
			19786: outdata = 32'd45750;
			19787: outdata = 32'd45749;
			19788: outdata = 32'd45748;
			19789: outdata = 32'd45747;
			19790: outdata = 32'd45746;
			19791: outdata = 32'd45745;
			19792: outdata = 32'd45744;
			19793: outdata = 32'd45743;
			19794: outdata = 32'd45742;
			19795: outdata = 32'd45741;
			19796: outdata = 32'd45740;
			19797: outdata = 32'd45739;
			19798: outdata = 32'd45738;
			19799: outdata = 32'd45737;
			19800: outdata = 32'd45736;
			19801: outdata = 32'd45735;
			19802: outdata = 32'd45734;
			19803: outdata = 32'd45733;
			19804: outdata = 32'd45732;
			19805: outdata = 32'd45731;
			19806: outdata = 32'd45730;
			19807: outdata = 32'd45729;
			19808: outdata = 32'd45728;
			19809: outdata = 32'd45727;
			19810: outdata = 32'd45726;
			19811: outdata = 32'd45725;
			19812: outdata = 32'd45724;
			19813: outdata = 32'd45723;
			19814: outdata = 32'd45722;
			19815: outdata = 32'd45721;
			19816: outdata = 32'd45720;
			19817: outdata = 32'd45719;
			19818: outdata = 32'd45718;
			19819: outdata = 32'd45717;
			19820: outdata = 32'd45716;
			19821: outdata = 32'd45715;
			19822: outdata = 32'd45714;
			19823: outdata = 32'd45713;
			19824: outdata = 32'd45712;
			19825: outdata = 32'd45711;
			19826: outdata = 32'd45710;
			19827: outdata = 32'd45709;
			19828: outdata = 32'd45708;
			19829: outdata = 32'd45707;
			19830: outdata = 32'd45706;
			19831: outdata = 32'd45705;
			19832: outdata = 32'd45704;
			19833: outdata = 32'd45703;
			19834: outdata = 32'd45702;
			19835: outdata = 32'd45701;
			19836: outdata = 32'd45700;
			19837: outdata = 32'd45699;
			19838: outdata = 32'd45698;
			19839: outdata = 32'd45697;
			19840: outdata = 32'd45696;
			19841: outdata = 32'd45695;
			19842: outdata = 32'd45694;
			19843: outdata = 32'd45693;
			19844: outdata = 32'd45692;
			19845: outdata = 32'd45691;
			19846: outdata = 32'd45690;
			19847: outdata = 32'd45689;
			19848: outdata = 32'd45688;
			19849: outdata = 32'd45687;
			19850: outdata = 32'd45686;
			19851: outdata = 32'd45685;
			19852: outdata = 32'd45684;
			19853: outdata = 32'd45683;
			19854: outdata = 32'd45682;
			19855: outdata = 32'd45681;
			19856: outdata = 32'd45680;
			19857: outdata = 32'd45679;
			19858: outdata = 32'd45678;
			19859: outdata = 32'd45677;
			19860: outdata = 32'd45676;
			19861: outdata = 32'd45675;
			19862: outdata = 32'd45674;
			19863: outdata = 32'd45673;
			19864: outdata = 32'd45672;
			19865: outdata = 32'd45671;
			19866: outdata = 32'd45670;
			19867: outdata = 32'd45669;
			19868: outdata = 32'd45668;
			19869: outdata = 32'd45667;
			19870: outdata = 32'd45666;
			19871: outdata = 32'd45665;
			19872: outdata = 32'd45664;
			19873: outdata = 32'd45663;
			19874: outdata = 32'd45662;
			19875: outdata = 32'd45661;
			19876: outdata = 32'd45660;
			19877: outdata = 32'd45659;
			19878: outdata = 32'd45658;
			19879: outdata = 32'd45657;
			19880: outdata = 32'd45656;
			19881: outdata = 32'd45655;
			19882: outdata = 32'd45654;
			19883: outdata = 32'd45653;
			19884: outdata = 32'd45652;
			19885: outdata = 32'd45651;
			19886: outdata = 32'd45650;
			19887: outdata = 32'd45649;
			19888: outdata = 32'd45648;
			19889: outdata = 32'd45647;
			19890: outdata = 32'd45646;
			19891: outdata = 32'd45645;
			19892: outdata = 32'd45644;
			19893: outdata = 32'd45643;
			19894: outdata = 32'd45642;
			19895: outdata = 32'd45641;
			19896: outdata = 32'd45640;
			19897: outdata = 32'd45639;
			19898: outdata = 32'd45638;
			19899: outdata = 32'd45637;
			19900: outdata = 32'd45636;
			19901: outdata = 32'd45635;
			19902: outdata = 32'd45634;
			19903: outdata = 32'd45633;
			19904: outdata = 32'd45632;
			19905: outdata = 32'd45631;
			19906: outdata = 32'd45630;
			19907: outdata = 32'd45629;
			19908: outdata = 32'd45628;
			19909: outdata = 32'd45627;
			19910: outdata = 32'd45626;
			19911: outdata = 32'd45625;
			19912: outdata = 32'd45624;
			19913: outdata = 32'd45623;
			19914: outdata = 32'd45622;
			19915: outdata = 32'd45621;
			19916: outdata = 32'd45620;
			19917: outdata = 32'd45619;
			19918: outdata = 32'd45618;
			19919: outdata = 32'd45617;
			19920: outdata = 32'd45616;
			19921: outdata = 32'd45615;
			19922: outdata = 32'd45614;
			19923: outdata = 32'd45613;
			19924: outdata = 32'd45612;
			19925: outdata = 32'd45611;
			19926: outdata = 32'd45610;
			19927: outdata = 32'd45609;
			19928: outdata = 32'd45608;
			19929: outdata = 32'd45607;
			19930: outdata = 32'd45606;
			19931: outdata = 32'd45605;
			19932: outdata = 32'd45604;
			19933: outdata = 32'd45603;
			19934: outdata = 32'd45602;
			19935: outdata = 32'd45601;
			19936: outdata = 32'd45600;
			19937: outdata = 32'd45599;
			19938: outdata = 32'd45598;
			19939: outdata = 32'd45597;
			19940: outdata = 32'd45596;
			19941: outdata = 32'd45595;
			19942: outdata = 32'd45594;
			19943: outdata = 32'd45593;
			19944: outdata = 32'd45592;
			19945: outdata = 32'd45591;
			19946: outdata = 32'd45590;
			19947: outdata = 32'd45589;
			19948: outdata = 32'd45588;
			19949: outdata = 32'd45587;
			19950: outdata = 32'd45586;
			19951: outdata = 32'd45585;
			19952: outdata = 32'd45584;
			19953: outdata = 32'd45583;
			19954: outdata = 32'd45582;
			19955: outdata = 32'd45581;
			19956: outdata = 32'd45580;
			19957: outdata = 32'd45579;
			19958: outdata = 32'd45578;
			19959: outdata = 32'd45577;
			19960: outdata = 32'd45576;
			19961: outdata = 32'd45575;
			19962: outdata = 32'd45574;
			19963: outdata = 32'd45573;
			19964: outdata = 32'd45572;
			19965: outdata = 32'd45571;
			19966: outdata = 32'd45570;
			19967: outdata = 32'd45569;
			19968: outdata = 32'd45568;
			19969: outdata = 32'd45567;
			19970: outdata = 32'd45566;
			19971: outdata = 32'd45565;
			19972: outdata = 32'd45564;
			19973: outdata = 32'd45563;
			19974: outdata = 32'd45562;
			19975: outdata = 32'd45561;
			19976: outdata = 32'd45560;
			19977: outdata = 32'd45559;
			19978: outdata = 32'd45558;
			19979: outdata = 32'd45557;
			19980: outdata = 32'd45556;
			19981: outdata = 32'd45555;
			19982: outdata = 32'd45554;
			19983: outdata = 32'd45553;
			19984: outdata = 32'd45552;
			19985: outdata = 32'd45551;
			19986: outdata = 32'd45550;
			19987: outdata = 32'd45549;
			19988: outdata = 32'd45548;
			19989: outdata = 32'd45547;
			19990: outdata = 32'd45546;
			19991: outdata = 32'd45545;
			19992: outdata = 32'd45544;
			19993: outdata = 32'd45543;
			19994: outdata = 32'd45542;
			19995: outdata = 32'd45541;
			19996: outdata = 32'd45540;
			19997: outdata = 32'd45539;
			19998: outdata = 32'd45538;
			19999: outdata = 32'd45537;
			20000: outdata = 32'd45536;
			20001: outdata = 32'd45535;
			20002: outdata = 32'd45534;
			20003: outdata = 32'd45533;
			20004: outdata = 32'd45532;
			20005: outdata = 32'd45531;
			20006: outdata = 32'd45530;
			20007: outdata = 32'd45529;
			20008: outdata = 32'd45528;
			20009: outdata = 32'd45527;
			20010: outdata = 32'd45526;
			20011: outdata = 32'd45525;
			20012: outdata = 32'd45524;
			20013: outdata = 32'd45523;
			20014: outdata = 32'd45522;
			20015: outdata = 32'd45521;
			20016: outdata = 32'd45520;
			20017: outdata = 32'd45519;
			20018: outdata = 32'd45518;
			20019: outdata = 32'd45517;
			20020: outdata = 32'd45516;
			20021: outdata = 32'd45515;
			20022: outdata = 32'd45514;
			20023: outdata = 32'd45513;
			20024: outdata = 32'd45512;
			20025: outdata = 32'd45511;
			20026: outdata = 32'd45510;
			20027: outdata = 32'd45509;
			20028: outdata = 32'd45508;
			20029: outdata = 32'd45507;
			20030: outdata = 32'd45506;
			20031: outdata = 32'd45505;
			20032: outdata = 32'd45504;
			20033: outdata = 32'd45503;
			20034: outdata = 32'd45502;
			20035: outdata = 32'd45501;
			20036: outdata = 32'd45500;
			20037: outdata = 32'd45499;
			20038: outdata = 32'd45498;
			20039: outdata = 32'd45497;
			20040: outdata = 32'd45496;
			20041: outdata = 32'd45495;
			20042: outdata = 32'd45494;
			20043: outdata = 32'd45493;
			20044: outdata = 32'd45492;
			20045: outdata = 32'd45491;
			20046: outdata = 32'd45490;
			20047: outdata = 32'd45489;
			20048: outdata = 32'd45488;
			20049: outdata = 32'd45487;
			20050: outdata = 32'd45486;
			20051: outdata = 32'd45485;
			20052: outdata = 32'd45484;
			20053: outdata = 32'd45483;
			20054: outdata = 32'd45482;
			20055: outdata = 32'd45481;
			20056: outdata = 32'd45480;
			20057: outdata = 32'd45479;
			20058: outdata = 32'd45478;
			20059: outdata = 32'd45477;
			20060: outdata = 32'd45476;
			20061: outdata = 32'd45475;
			20062: outdata = 32'd45474;
			20063: outdata = 32'd45473;
			20064: outdata = 32'd45472;
			20065: outdata = 32'd45471;
			20066: outdata = 32'd45470;
			20067: outdata = 32'd45469;
			20068: outdata = 32'd45468;
			20069: outdata = 32'd45467;
			20070: outdata = 32'd45466;
			20071: outdata = 32'd45465;
			20072: outdata = 32'd45464;
			20073: outdata = 32'd45463;
			20074: outdata = 32'd45462;
			20075: outdata = 32'd45461;
			20076: outdata = 32'd45460;
			20077: outdata = 32'd45459;
			20078: outdata = 32'd45458;
			20079: outdata = 32'd45457;
			20080: outdata = 32'd45456;
			20081: outdata = 32'd45455;
			20082: outdata = 32'd45454;
			20083: outdata = 32'd45453;
			20084: outdata = 32'd45452;
			20085: outdata = 32'd45451;
			20086: outdata = 32'd45450;
			20087: outdata = 32'd45449;
			20088: outdata = 32'd45448;
			20089: outdata = 32'd45447;
			20090: outdata = 32'd45446;
			20091: outdata = 32'd45445;
			20092: outdata = 32'd45444;
			20093: outdata = 32'd45443;
			20094: outdata = 32'd45442;
			20095: outdata = 32'd45441;
			20096: outdata = 32'd45440;
			20097: outdata = 32'd45439;
			20098: outdata = 32'd45438;
			20099: outdata = 32'd45437;
			20100: outdata = 32'd45436;
			20101: outdata = 32'd45435;
			20102: outdata = 32'd45434;
			20103: outdata = 32'd45433;
			20104: outdata = 32'd45432;
			20105: outdata = 32'd45431;
			20106: outdata = 32'd45430;
			20107: outdata = 32'd45429;
			20108: outdata = 32'd45428;
			20109: outdata = 32'd45427;
			20110: outdata = 32'd45426;
			20111: outdata = 32'd45425;
			20112: outdata = 32'd45424;
			20113: outdata = 32'd45423;
			20114: outdata = 32'd45422;
			20115: outdata = 32'd45421;
			20116: outdata = 32'd45420;
			20117: outdata = 32'd45419;
			20118: outdata = 32'd45418;
			20119: outdata = 32'd45417;
			20120: outdata = 32'd45416;
			20121: outdata = 32'd45415;
			20122: outdata = 32'd45414;
			20123: outdata = 32'd45413;
			20124: outdata = 32'd45412;
			20125: outdata = 32'd45411;
			20126: outdata = 32'd45410;
			20127: outdata = 32'd45409;
			20128: outdata = 32'd45408;
			20129: outdata = 32'd45407;
			20130: outdata = 32'd45406;
			20131: outdata = 32'd45405;
			20132: outdata = 32'd45404;
			20133: outdata = 32'd45403;
			20134: outdata = 32'd45402;
			20135: outdata = 32'd45401;
			20136: outdata = 32'd45400;
			20137: outdata = 32'd45399;
			20138: outdata = 32'd45398;
			20139: outdata = 32'd45397;
			20140: outdata = 32'd45396;
			20141: outdata = 32'd45395;
			20142: outdata = 32'd45394;
			20143: outdata = 32'd45393;
			20144: outdata = 32'd45392;
			20145: outdata = 32'd45391;
			20146: outdata = 32'd45390;
			20147: outdata = 32'd45389;
			20148: outdata = 32'd45388;
			20149: outdata = 32'd45387;
			20150: outdata = 32'd45386;
			20151: outdata = 32'd45385;
			20152: outdata = 32'd45384;
			20153: outdata = 32'd45383;
			20154: outdata = 32'd45382;
			20155: outdata = 32'd45381;
			20156: outdata = 32'd45380;
			20157: outdata = 32'd45379;
			20158: outdata = 32'd45378;
			20159: outdata = 32'd45377;
			20160: outdata = 32'd45376;
			20161: outdata = 32'd45375;
			20162: outdata = 32'd45374;
			20163: outdata = 32'd45373;
			20164: outdata = 32'd45372;
			20165: outdata = 32'd45371;
			20166: outdata = 32'd45370;
			20167: outdata = 32'd45369;
			20168: outdata = 32'd45368;
			20169: outdata = 32'd45367;
			20170: outdata = 32'd45366;
			20171: outdata = 32'd45365;
			20172: outdata = 32'd45364;
			20173: outdata = 32'd45363;
			20174: outdata = 32'd45362;
			20175: outdata = 32'd45361;
			20176: outdata = 32'd45360;
			20177: outdata = 32'd45359;
			20178: outdata = 32'd45358;
			20179: outdata = 32'd45357;
			20180: outdata = 32'd45356;
			20181: outdata = 32'd45355;
			20182: outdata = 32'd45354;
			20183: outdata = 32'd45353;
			20184: outdata = 32'd45352;
			20185: outdata = 32'd45351;
			20186: outdata = 32'd45350;
			20187: outdata = 32'd45349;
			20188: outdata = 32'd45348;
			20189: outdata = 32'd45347;
			20190: outdata = 32'd45346;
			20191: outdata = 32'd45345;
			20192: outdata = 32'd45344;
			20193: outdata = 32'd45343;
			20194: outdata = 32'd45342;
			20195: outdata = 32'd45341;
			20196: outdata = 32'd45340;
			20197: outdata = 32'd45339;
			20198: outdata = 32'd45338;
			20199: outdata = 32'd45337;
			20200: outdata = 32'd45336;
			20201: outdata = 32'd45335;
			20202: outdata = 32'd45334;
			20203: outdata = 32'd45333;
			20204: outdata = 32'd45332;
			20205: outdata = 32'd45331;
			20206: outdata = 32'd45330;
			20207: outdata = 32'd45329;
			20208: outdata = 32'd45328;
			20209: outdata = 32'd45327;
			20210: outdata = 32'd45326;
			20211: outdata = 32'd45325;
			20212: outdata = 32'd45324;
			20213: outdata = 32'd45323;
			20214: outdata = 32'd45322;
			20215: outdata = 32'd45321;
			20216: outdata = 32'd45320;
			20217: outdata = 32'd45319;
			20218: outdata = 32'd45318;
			20219: outdata = 32'd45317;
			20220: outdata = 32'd45316;
			20221: outdata = 32'd45315;
			20222: outdata = 32'd45314;
			20223: outdata = 32'd45313;
			20224: outdata = 32'd45312;
			20225: outdata = 32'd45311;
			20226: outdata = 32'd45310;
			20227: outdata = 32'd45309;
			20228: outdata = 32'd45308;
			20229: outdata = 32'd45307;
			20230: outdata = 32'd45306;
			20231: outdata = 32'd45305;
			20232: outdata = 32'd45304;
			20233: outdata = 32'd45303;
			20234: outdata = 32'd45302;
			20235: outdata = 32'd45301;
			20236: outdata = 32'd45300;
			20237: outdata = 32'd45299;
			20238: outdata = 32'd45298;
			20239: outdata = 32'd45297;
			20240: outdata = 32'd45296;
			20241: outdata = 32'd45295;
			20242: outdata = 32'd45294;
			20243: outdata = 32'd45293;
			20244: outdata = 32'd45292;
			20245: outdata = 32'd45291;
			20246: outdata = 32'd45290;
			20247: outdata = 32'd45289;
			20248: outdata = 32'd45288;
			20249: outdata = 32'd45287;
			20250: outdata = 32'd45286;
			20251: outdata = 32'd45285;
			20252: outdata = 32'd45284;
			20253: outdata = 32'd45283;
			20254: outdata = 32'd45282;
			20255: outdata = 32'd45281;
			20256: outdata = 32'd45280;
			20257: outdata = 32'd45279;
			20258: outdata = 32'd45278;
			20259: outdata = 32'd45277;
			20260: outdata = 32'd45276;
			20261: outdata = 32'd45275;
			20262: outdata = 32'd45274;
			20263: outdata = 32'd45273;
			20264: outdata = 32'd45272;
			20265: outdata = 32'd45271;
			20266: outdata = 32'd45270;
			20267: outdata = 32'd45269;
			20268: outdata = 32'd45268;
			20269: outdata = 32'd45267;
			20270: outdata = 32'd45266;
			20271: outdata = 32'd45265;
			20272: outdata = 32'd45264;
			20273: outdata = 32'd45263;
			20274: outdata = 32'd45262;
			20275: outdata = 32'd45261;
			20276: outdata = 32'd45260;
			20277: outdata = 32'd45259;
			20278: outdata = 32'd45258;
			20279: outdata = 32'd45257;
			20280: outdata = 32'd45256;
			20281: outdata = 32'd45255;
			20282: outdata = 32'd45254;
			20283: outdata = 32'd45253;
			20284: outdata = 32'd45252;
			20285: outdata = 32'd45251;
			20286: outdata = 32'd45250;
			20287: outdata = 32'd45249;
			20288: outdata = 32'd45248;
			20289: outdata = 32'd45247;
			20290: outdata = 32'd45246;
			20291: outdata = 32'd45245;
			20292: outdata = 32'd45244;
			20293: outdata = 32'd45243;
			20294: outdata = 32'd45242;
			20295: outdata = 32'd45241;
			20296: outdata = 32'd45240;
			20297: outdata = 32'd45239;
			20298: outdata = 32'd45238;
			20299: outdata = 32'd45237;
			20300: outdata = 32'd45236;
			20301: outdata = 32'd45235;
			20302: outdata = 32'd45234;
			20303: outdata = 32'd45233;
			20304: outdata = 32'd45232;
			20305: outdata = 32'd45231;
			20306: outdata = 32'd45230;
			20307: outdata = 32'd45229;
			20308: outdata = 32'd45228;
			20309: outdata = 32'd45227;
			20310: outdata = 32'd45226;
			20311: outdata = 32'd45225;
			20312: outdata = 32'd45224;
			20313: outdata = 32'd45223;
			20314: outdata = 32'd45222;
			20315: outdata = 32'd45221;
			20316: outdata = 32'd45220;
			20317: outdata = 32'd45219;
			20318: outdata = 32'd45218;
			20319: outdata = 32'd45217;
			20320: outdata = 32'd45216;
			20321: outdata = 32'd45215;
			20322: outdata = 32'd45214;
			20323: outdata = 32'd45213;
			20324: outdata = 32'd45212;
			20325: outdata = 32'd45211;
			20326: outdata = 32'd45210;
			20327: outdata = 32'd45209;
			20328: outdata = 32'd45208;
			20329: outdata = 32'd45207;
			20330: outdata = 32'd45206;
			20331: outdata = 32'd45205;
			20332: outdata = 32'd45204;
			20333: outdata = 32'd45203;
			20334: outdata = 32'd45202;
			20335: outdata = 32'd45201;
			20336: outdata = 32'd45200;
			20337: outdata = 32'd45199;
			20338: outdata = 32'd45198;
			20339: outdata = 32'd45197;
			20340: outdata = 32'd45196;
			20341: outdata = 32'd45195;
			20342: outdata = 32'd45194;
			20343: outdata = 32'd45193;
			20344: outdata = 32'd45192;
			20345: outdata = 32'd45191;
			20346: outdata = 32'd45190;
			20347: outdata = 32'd45189;
			20348: outdata = 32'd45188;
			20349: outdata = 32'd45187;
			20350: outdata = 32'd45186;
			20351: outdata = 32'd45185;
			20352: outdata = 32'd45184;
			20353: outdata = 32'd45183;
			20354: outdata = 32'd45182;
			20355: outdata = 32'd45181;
			20356: outdata = 32'd45180;
			20357: outdata = 32'd45179;
			20358: outdata = 32'd45178;
			20359: outdata = 32'd45177;
			20360: outdata = 32'd45176;
			20361: outdata = 32'd45175;
			20362: outdata = 32'd45174;
			20363: outdata = 32'd45173;
			20364: outdata = 32'd45172;
			20365: outdata = 32'd45171;
			20366: outdata = 32'd45170;
			20367: outdata = 32'd45169;
			20368: outdata = 32'd45168;
			20369: outdata = 32'd45167;
			20370: outdata = 32'd45166;
			20371: outdata = 32'd45165;
			20372: outdata = 32'd45164;
			20373: outdata = 32'd45163;
			20374: outdata = 32'd45162;
			20375: outdata = 32'd45161;
			20376: outdata = 32'd45160;
			20377: outdata = 32'd45159;
			20378: outdata = 32'd45158;
			20379: outdata = 32'd45157;
			20380: outdata = 32'd45156;
			20381: outdata = 32'd45155;
			20382: outdata = 32'd45154;
			20383: outdata = 32'd45153;
			20384: outdata = 32'd45152;
			20385: outdata = 32'd45151;
			20386: outdata = 32'd45150;
			20387: outdata = 32'd45149;
			20388: outdata = 32'd45148;
			20389: outdata = 32'd45147;
			20390: outdata = 32'd45146;
			20391: outdata = 32'd45145;
			20392: outdata = 32'd45144;
			20393: outdata = 32'd45143;
			20394: outdata = 32'd45142;
			20395: outdata = 32'd45141;
			20396: outdata = 32'd45140;
			20397: outdata = 32'd45139;
			20398: outdata = 32'd45138;
			20399: outdata = 32'd45137;
			20400: outdata = 32'd45136;
			20401: outdata = 32'd45135;
			20402: outdata = 32'd45134;
			20403: outdata = 32'd45133;
			20404: outdata = 32'd45132;
			20405: outdata = 32'd45131;
			20406: outdata = 32'd45130;
			20407: outdata = 32'd45129;
			20408: outdata = 32'd45128;
			20409: outdata = 32'd45127;
			20410: outdata = 32'd45126;
			20411: outdata = 32'd45125;
			20412: outdata = 32'd45124;
			20413: outdata = 32'd45123;
			20414: outdata = 32'd45122;
			20415: outdata = 32'd45121;
			20416: outdata = 32'd45120;
			20417: outdata = 32'd45119;
			20418: outdata = 32'd45118;
			20419: outdata = 32'd45117;
			20420: outdata = 32'd45116;
			20421: outdata = 32'd45115;
			20422: outdata = 32'd45114;
			20423: outdata = 32'd45113;
			20424: outdata = 32'd45112;
			20425: outdata = 32'd45111;
			20426: outdata = 32'd45110;
			20427: outdata = 32'd45109;
			20428: outdata = 32'd45108;
			20429: outdata = 32'd45107;
			20430: outdata = 32'd45106;
			20431: outdata = 32'd45105;
			20432: outdata = 32'd45104;
			20433: outdata = 32'd45103;
			20434: outdata = 32'd45102;
			20435: outdata = 32'd45101;
			20436: outdata = 32'd45100;
			20437: outdata = 32'd45099;
			20438: outdata = 32'd45098;
			20439: outdata = 32'd45097;
			20440: outdata = 32'd45096;
			20441: outdata = 32'd45095;
			20442: outdata = 32'd45094;
			20443: outdata = 32'd45093;
			20444: outdata = 32'd45092;
			20445: outdata = 32'd45091;
			20446: outdata = 32'd45090;
			20447: outdata = 32'd45089;
			20448: outdata = 32'd45088;
			20449: outdata = 32'd45087;
			20450: outdata = 32'd45086;
			20451: outdata = 32'd45085;
			20452: outdata = 32'd45084;
			20453: outdata = 32'd45083;
			20454: outdata = 32'd45082;
			20455: outdata = 32'd45081;
			20456: outdata = 32'd45080;
			20457: outdata = 32'd45079;
			20458: outdata = 32'd45078;
			20459: outdata = 32'd45077;
			20460: outdata = 32'd45076;
			20461: outdata = 32'd45075;
			20462: outdata = 32'd45074;
			20463: outdata = 32'd45073;
			20464: outdata = 32'd45072;
			20465: outdata = 32'd45071;
			20466: outdata = 32'd45070;
			20467: outdata = 32'd45069;
			20468: outdata = 32'd45068;
			20469: outdata = 32'd45067;
			20470: outdata = 32'd45066;
			20471: outdata = 32'd45065;
			20472: outdata = 32'd45064;
			20473: outdata = 32'd45063;
			20474: outdata = 32'd45062;
			20475: outdata = 32'd45061;
			20476: outdata = 32'd45060;
			20477: outdata = 32'd45059;
			20478: outdata = 32'd45058;
			20479: outdata = 32'd45057;
			20480: outdata = 32'd45056;
			20481: outdata = 32'd45055;
			20482: outdata = 32'd45054;
			20483: outdata = 32'd45053;
			20484: outdata = 32'd45052;
			20485: outdata = 32'd45051;
			20486: outdata = 32'd45050;
			20487: outdata = 32'd45049;
			20488: outdata = 32'd45048;
			20489: outdata = 32'd45047;
			20490: outdata = 32'd45046;
			20491: outdata = 32'd45045;
			20492: outdata = 32'd45044;
			20493: outdata = 32'd45043;
			20494: outdata = 32'd45042;
			20495: outdata = 32'd45041;
			20496: outdata = 32'd45040;
			20497: outdata = 32'd45039;
			20498: outdata = 32'd45038;
			20499: outdata = 32'd45037;
			20500: outdata = 32'd45036;
			20501: outdata = 32'd45035;
			20502: outdata = 32'd45034;
			20503: outdata = 32'd45033;
			20504: outdata = 32'd45032;
			20505: outdata = 32'd45031;
			20506: outdata = 32'd45030;
			20507: outdata = 32'd45029;
			20508: outdata = 32'd45028;
			20509: outdata = 32'd45027;
			20510: outdata = 32'd45026;
			20511: outdata = 32'd45025;
			20512: outdata = 32'd45024;
			20513: outdata = 32'd45023;
			20514: outdata = 32'd45022;
			20515: outdata = 32'd45021;
			20516: outdata = 32'd45020;
			20517: outdata = 32'd45019;
			20518: outdata = 32'd45018;
			20519: outdata = 32'd45017;
			20520: outdata = 32'd45016;
			20521: outdata = 32'd45015;
			20522: outdata = 32'd45014;
			20523: outdata = 32'd45013;
			20524: outdata = 32'd45012;
			20525: outdata = 32'd45011;
			20526: outdata = 32'd45010;
			20527: outdata = 32'd45009;
			20528: outdata = 32'd45008;
			20529: outdata = 32'd45007;
			20530: outdata = 32'd45006;
			20531: outdata = 32'd45005;
			20532: outdata = 32'd45004;
			20533: outdata = 32'd45003;
			20534: outdata = 32'd45002;
			20535: outdata = 32'd45001;
			20536: outdata = 32'd45000;
			20537: outdata = 32'd44999;
			20538: outdata = 32'd44998;
			20539: outdata = 32'd44997;
			20540: outdata = 32'd44996;
			20541: outdata = 32'd44995;
			20542: outdata = 32'd44994;
			20543: outdata = 32'd44993;
			20544: outdata = 32'd44992;
			20545: outdata = 32'd44991;
			20546: outdata = 32'd44990;
			20547: outdata = 32'd44989;
			20548: outdata = 32'd44988;
			20549: outdata = 32'd44987;
			20550: outdata = 32'd44986;
			20551: outdata = 32'd44985;
			20552: outdata = 32'd44984;
			20553: outdata = 32'd44983;
			20554: outdata = 32'd44982;
			20555: outdata = 32'd44981;
			20556: outdata = 32'd44980;
			20557: outdata = 32'd44979;
			20558: outdata = 32'd44978;
			20559: outdata = 32'd44977;
			20560: outdata = 32'd44976;
			20561: outdata = 32'd44975;
			20562: outdata = 32'd44974;
			20563: outdata = 32'd44973;
			20564: outdata = 32'd44972;
			20565: outdata = 32'd44971;
			20566: outdata = 32'd44970;
			20567: outdata = 32'd44969;
			20568: outdata = 32'd44968;
			20569: outdata = 32'd44967;
			20570: outdata = 32'd44966;
			20571: outdata = 32'd44965;
			20572: outdata = 32'd44964;
			20573: outdata = 32'd44963;
			20574: outdata = 32'd44962;
			20575: outdata = 32'd44961;
			20576: outdata = 32'd44960;
			20577: outdata = 32'd44959;
			20578: outdata = 32'd44958;
			20579: outdata = 32'd44957;
			20580: outdata = 32'd44956;
			20581: outdata = 32'd44955;
			20582: outdata = 32'd44954;
			20583: outdata = 32'd44953;
			20584: outdata = 32'd44952;
			20585: outdata = 32'd44951;
			20586: outdata = 32'd44950;
			20587: outdata = 32'd44949;
			20588: outdata = 32'd44948;
			20589: outdata = 32'd44947;
			20590: outdata = 32'd44946;
			20591: outdata = 32'd44945;
			20592: outdata = 32'd44944;
			20593: outdata = 32'd44943;
			20594: outdata = 32'd44942;
			20595: outdata = 32'd44941;
			20596: outdata = 32'd44940;
			20597: outdata = 32'd44939;
			20598: outdata = 32'd44938;
			20599: outdata = 32'd44937;
			20600: outdata = 32'd44936;
			20601: outdata = 32'd44935;
			20602: outdata = 32'd44934;
			20603: outdata = 32'd44933;
			20604: outdata = 32'd44932;
			20605: outdata = 32'd44931;
			20606: outdata = 32'd44930;
			20607: outdata = 32'd44929;
			20608: outdata = 32'd44928;
			20609: outdata = 32'd44927;
			20610: outdata = 32'd44926;
			20611: outdata = 32'd44925;
			20612: outdata = 32'd44924;
			20613: outdata = 32'd44923;
			20614: outdata = 32'd44922;
			20615: outdata = 32'd44921;
			20616: outdata = 32'd44920;
			20617: outdata = 32'd44919;
			20618: outdata = 32'd44918;
			20619: outdata = 32'd44917;
			20620: outdata = 32'd44916;
			20621: outdata = 32'd44915;
			20622: outdata = 32'd44914;
			20623: outdata = 32'd44913;
			20624: outdata = 32'd44912;
			20625: outdata = 32'd44911;
			20626: outdata = 32'd44910;
			20627: outdata = 32'd44909;
			20628: outdata = 32'd44908;
			20629: outdata = 32'd44907;
			20630: outdata = 32'd44906;
			20631: outdata = 32'd44905;
			20632: outdata = 32'd44904;
			20633: outdata = 32'd44903;
			20634: outdata = 32'd44902;
			20635: outdata = 32'd44901;
			20636: outdata = 32'd44900;
			20637: outdata = 32'd44899;
			20638: outdata = 32'd44898;
			20639: outdata = 32'd44897;
			20640: outdata = 32'd44896;
			20641: outdata = 32'd44895;
			20642: outdata = 32'd44894;
			20643: outdata = 32'd44893;
			20644: outdata = 32'd44892;
			20645: outdata = 32'd44891;
			20646: outdata = 32'd44890;
			20647: outdata = 32'd44889;
			20648: outdata = 32'd44888;
			20649: outdata = 32'd44887;
			20650: outdata = 32'd44886;
			20651: outdata = 32'd44885;
			20652: outdata = 32'd44884;
			20653: outdata = 32'd44883;
			20654: outdata = 32'd44882;
			20655: outdata = 32'd44881;
			20656: outdata = 32'd44880;
			20657: outdata = 32'd44879;
			20658: outdata = 32'd44878;
			20659: outdata = 32'd44877;
			20660: outdata = 32'd44876;
			20661: outdata = 32'd44875;
			20662: outdata = 32'd44874;
			20663: outdata = 32'd44873;
			20664: outdata = 32'd44872;
			20665: outdata = 32'd44871;
			20666: outdata = 32'd44870;
			20667: outdata = 32'd44869;
			20668: outdata = 32'd44868;
			20669: outdata = 32'd44867;
			20670: outdata = 32'd44866;
			20671: outdata = 32'd44865;
			20672: outdata = 32'd44864;
			20673: outdata = 32'd44863;
			20674: outdata = 32'd44862;
			20675: outdata = 32'd44861;
			20676: outdata = 32'd44860;
			20677: outdata = 32'd44859;
			20678: outdata = 32'd44858;
			20679: outdata = 32'd44857;
			20680: outdata = 32'd44856;
			20681: outdata = 32'd44855;
			20682: outdata = 32'd44854;
			20683: outdata = 32'd44853;
			20684: outdata = 32'd44852;
			20685: outdata = 32'd44851;
			20686: outdata = 32'd44850;
			20687: outdata = 32'd44849;
			20688: outdata = 32'd44848;
			20689: outdata = 32'd44847;
			20690: outdata = 32'd44846;
			20691: outdata = 32'd44845;
			20692: outdata = 32'd44844;
			20693: outdata = 32'd44843;
			20694: outdata = 32'd44842;
			20695: outdata = 32'd44841;
			20696: outdata = 32'd44840;
			20697: outdata = 32'd44839;
			20698: outdata = 32'd44838;
			20699: outdata = 32'd44837;
			20700: outdata = 32'd44836;
			20701: outdata = 32'd44835;
			20702: outdata = 32'd44834;
			20703: outdata = 32'd44833;
			20704: outdata = 32'd44832;
			20705: outdata = 32'd44831;
			20706: outdata = 32'd44830;
			20707: outdata = 32'd44829;
			20708: outdata = 32'd44828;
			20709: outdata = 32'd44827;
			20710: outdata = 32'd44826;
			20711: outdata = 32'd44825;
			20712: outdata = 32'd44824;
			20713: outdata = 32'd44823;
			20714: outdata = 32'd44822;
			20715: outdata = 32'd44821;
			20716: outdata = 32'd44820;
			20717: outdata = 32'd44819;
			20718: outdata = 32'd44818;
			20719: outdata = 32'd44817;
			20720: outdata = 32'd44816;
			20721: outdata = 32'd44815;
			20722: outdata = 32'd44814;
			20723: outdata = 32'd44813;
			20724: outdata = 32'd44812;
			20725: outdata = 32'd44811;
			20726: outdata = 32'd44810;
			20727: outdata = 32'd44809;
			20728: outdata = 32'd44808;
			20729: outdata = 32'd44807;
			20730: outdata = 32'd44806;
			20731: outdata = 32'd44805;
			20732: outdata = 32'd44804;
			20733: outdata = 32'd44803;
			20734: outdata = 32'd44802;
			20735: outdata = 32'd44801;
			20736: outdata = 32'd44800;
			20737: outdata = 32'd44799;
			20738: outdata = 32'd44798;
			20739: outdata = 32'd44797;
			20740: outdata = 32'd44796;
			20741: outdata = 32'd44795;
			20742: outdata = 32'd44794;
			20743: outdata = 32'd44793;
			20744: outdata = 32'd44792;
			20745: outdata = 32'd44791;
			20746: outdata = 32'd44790;
			20747: outdata = 32'd44789;
			20748: outdata = 32'd44788;
			20749: outdata = 32'd44787;
			20750: outdata = 32'd44786;
			20751: outdata = 32'd44785;
			20752: outdata = 32'd44784;
			20753: outdata = 32'd44783;
			20754: outdata = 32'd44782;
			20755: outdata = 32'd44781;
			20756: outdata = 32'd44780;
			20757: outdata = 32'd44779;
			20758: outdata = 32'd44778;
			20759: outdata = 32'd44777;
			20760: outdata = 32'd44776;
			20761: outdata = 32'd44775;
			20762: outdata = 32'd44774;
			20763: outdata = 32'd44773;
			20764: outdata = 32'd44772;
			20765: outdata = 32'd44771;
			20766: outdata = 32'd44770;
			20767: outdata = 32'd44769;
			20768: outdata = 32'd44768;
			20769: outdata = 32'd44767;
			20770: outdata = 32'd44766;
			20771: outdata = 32'd44765;
			20772: outdata = 32'd44764;
			20773: outdata = 32'd44763;
			20774: outdata = 32'd44762;
			20775: outdata = 32'd44761;
			20776: outdata = 32'd44760;
			20777: outdata = 32'd44759;
			20778: outdata = 32'd44758;
			20779: outdata = 32'd44757;
			20780: outdata = 32'd44756;
			20781: outdata = 32'd44755;
			20782: outdata = 32'd44754;
			20783: outdata = 32'd44753;
			20784: outdata = 32'd44752;
			20785: outdata = 32'd44751;
			20786: outdata = 32'd44750;
			20787: outdata = 32'd44749;
			20788: outdata = 32'd44748;
			20789: outdata = 32'd44747;
			20790: outdata = 32'd44746;
			20791: outdata = 32'd44745;
			20792: outdata = 32'd44744;
			20793: outdata = 32'd44743;
			20794: outdata = 32'd44742;
			20795: outdata = 32'd44741;
			20796: outdata = 32'd44740;
			20797: outdata = 32'd44739;
			20798: outdata = 32'd44738;
			20799: outdata = 32'd44737;
			20800: outdata = 32'd44736;
			20801: outdata = 32'd44735;
			20802: outdata = 32'd44734;
			20803: outdata = 32'd44733;
			20804: outdata = 32'd44732;
			20805: outdata = 32'd44731;
			20806: outdata = 32'd44730;
			20807: outdata = 32'd44729;
			20808: outdata = 32'd44728;
			20809: outdata = 32'd44727;
			20810: outdata = 32'd44726;
			20811: outdata = 32'd44725;
			20812: outdata = 32'd44724;
			20813: outdata = 32'd44723;
			20814: outdata = 32'd44722;
			20815: outdata = 32'd44721;
			20816: outdata = 32'd44720;
			20817: outdata = 32'd44719;
			20818: outdata = 32'd44718;
			20819: outdata = 32'd44717;
			20820: outdata = 32'd44716;
			20821: outdata = 32'd44715;
			20822: outdata = 32'd44714;
			20823: outdata = 32'd44713;
			20824: outdata = 32'd44712;
			20825: outdata = 32'd44711;
			20826: outdata = 32'd44710;
			20827: outdata = 32'd44709;
			20828: outdata = 32'd44708;
			20829: outdata = 32'd44707;
			20830: outdata = 32'd44706;
			20831: outdata = 32'd44705;
			20832: outdata = 32'd44704;
			20833: outdata = 32'd44703;
			20834: outdata = 32'd44702;
			20835: outdata = 32'd44701;
			20836: outdata = 32'd44700;
			20837: outdata = 32'd44699;
			20838: outdata = 32'd44698;
			20839: outdata = 32'd44697;
			20840: outdata = 32'd44696;
			20841: outdata = 32'd44695;
			20842: outdata = 32'd44694;
			20843: outdata = 32'd44693;
			20844: outdata = 32'd44692;
			20845: outdata = 32'd44691;
			20846: outdata = 32'd44690;
			20847: outdata = 32'd44689;
			20848: outdata = 32'd44688;
			20849: outdata = 32'd44687;
			20850: outdata = 32'd44686;
			20851: outdata = 32'd44685;
			20852: outdata = 32'd44684;
			20853: outdata = 32'd44683;
			20854: outdata = 32'd44682;
			20855: outdata = 32'd44681;
			20856: outdata = 32'd44680;
			20857: outdata = 32'd44679;
			20858: outdata = 32'd44678;
			20859: outdata = 32'd44677;
			20860: outdata = 32'd44676;
			20861: outdata = 32'd44675;
			20862: outdata = 32'd44674;
			20863: outdata = 32'd44673;
			20864: outdata = 32'd44672;
			20865: outdata = 32'd44671;
			20866: outdata = 32'd44670;
			20867: outdata = 32'd44669;
			20868: outdata = 32'd44668;
			20869: outdata = 32'd44667;
			20870: outdata = 32'd44666;
			20871: outdata = 32'd44665;
			20872: outdata = 32'd44664;
			20873: outdata = 32'd44663;
			20874: outdata = 32'd44662;
			20875: outdata = 32'd44661;
			20876: outdata = 32'd44660;
			20877: outdata = 32'd44659;
			20878: outdata = 32'd44658;
			20879: outdata = 32'd44657;
			20880: outdata = 32'd44656;
			20881: outdata = 32'd44655;
			20882: outdata = 32'd44654;
			20883: outdata = 32'd44653;
			20884: outdata = 32'd44652;
			20885: outdata = 32'd44651;
			20886: outdata = 32'd44650;
			20887: outdata = 32'd44649;
			20888: outdata = 32'd44648;
			20889: outdata = 32'd44647;
			20890: outdata = 32'd44646;
			20891: outdata = 32'd44645;
			20892: outdata = 32'd44644;
			20893: outdata = 32'd44643;
			20894: outdata = 32'd44642;
			20895: outdata = 32'd44641;
			20896: outdata = 32'd44640;
			20897: outdata = 32'd44639;
			20898: outdata = 32'd44638;
			20899: outdata = 32'd44637;
			20900: outdata = 32'd44636;
			20901: outdata = 32'd44635;
			20902: outdata = 32'd44634;
			20903: outdata = 32'd44633;
			20904: outdata = 32'd44632;
			20905: outdata = 32'd44631;
			20906: outdata = 32'd44630;
			20907: outdata = 32'd44629;
			20908: outdata = 32'd44628;
			20909: outdata = 32'd44627;
			20910: outdata = 32'd44626;
			20911: outdata = 32'd44625;
			20912: outdata = 32'd44624;
			20913: outdata = 32'd44623;
			20914: outdata = 32'd44622;
			20915: outdata = 32'd44621;
			20916: outdata = 32'd44620;
			20917: outdata = 32'd44619;
			20918: outdata = 32'd44618;
			20919: outdata = 32'd44617;
			20920: outdata = 32'd44616;
			20921: outdata = 32'd44615;
			20922: outdata = 32'd44614;
			20923: outdata = 32'd44613;
			20924: outdata = 32'd44612;
			20925: outdata = 32'd44611;
			20926: outdata = 32'd44610;
			20927: outdata = 32'd44609;
			20928: outdata = 32'd44608;
			20929: outdata = 32'd44607;
			20930: outdata = 32'd44606;
			20931: outdata = 32'd44605;
			20932: outdata = 32'd44604;
			20933: outdata = 32'd44603;
			20934: outdata = 32'd44602;
			20935: outdata = 32'd44601;
			20936: outdata = 32'd44600;
			20937: outdata = 32'd44599;
			20938: outdata = 32'd44598;
			20939: outdata = 32'd44597;
			20940: outdata = 32'd44596;
			20941: outdata = 32'd44595;
			20942: outdata = 32'd44594;
			20943: outdata = 32'd44593;
			20944: outdata = 32'd44592;
			20945: outdata = 32'd44591;
			20946: outdata = 32'd44590;
			20947: outdata = 32'd44589;
			20948: outdata = 32'd44588;
			20949: outdata = 32'd44587;
			20950: outdata = 32'd44586;
			20951: outdata = 32'd44585;
			20952: outdata = 32'd44584;
			20953: outdata = 32'd44583;
			20954: outdata = 32'd44582;
			20955: outdata = 32'd44581;
			20956: outdata = 32'd44580;
			20957: outdata = 32'd44579;
			20958: outdata = 32'd44578;
			20959: outdata = 32'd44577;
			20960: outdata = 32'd44576;
			20961: outdata = 32'd44575;
			20962: outdata = 32'd44574;
			20963: outdata = 32'd44573;
			20964: outdata = 32'd44572;
			20965: outdata = 32'd44571;
			20966: outdata = 32'd44570;
			20967: outdata = 32'd44569;
			20968: outdata = 32'd44568;
			20969: outdata = 32'd44567;
			20970: outdata = 32'd44566;
			20971: outdata = 32'd44565;
			20972: outdata = 32'd44564;
			20973: outdata = 32'd44563;
			20974: outdata = 32'd44562;
			20975: outdata = 32'd44561;
			20976: outdata = 32'd44560;
			20977: outdata = 32'd44559;
			20978: outdata = 32'd44558;
			20979: outdata = 32'd44557;
			20980: outdata = 32'd44556;
			20981: outdata = 32'd44555;
			20982: outdata = 32'd44554;
			20983: outdata = 32'd44553;
			20984: outdata = 32'd44552;
			20985: outdata = 32'd44551;
			20986: outdata = 32'd44550;
			20987: outdata = 32'd44549;
			20988: outdata = 32'd44548;
			20989: outdata = 32'd44547;
			20990: outdata = 32'd44546;
			20991: outdata = 32'd44545;
			20992: outdata = 32'd44544;
			20993: outdata = 32'd44543;
			20994: outdata = 32'd44542;
			20995: outdata = 32'd44541;
			20996: outdata = 32'd44540;
			20997: outdata = 32'd44539;
			20998: outdata = 32'd44538;
			20999: outdata = 32'd44537;
			21000: outdata = 32'd44536;
			21001: outdata = 32'd44535;
			21002: outdata = 32'd44534;
			21003: outdata = 32'd44533;
			21004: outdata = 32'd44532;
			21005: outdata = 32'd44531;
			21006: outdata = 32'd44530;
			21007: outdata = 32'd44529;
			21008: outdata = 32'd44528;
			21009: outdata = 32'd44527;
			21010: outdata = 32'd44526;
			21011: outdata = 32'd44525;
			21012: outdata = 32'd44524;
			21013: outdata = 32'd44523;
			21014: outdata = 32'd44522;
			21015: outdata = 32'd44521;
			21016: outdata = 32'd44520;
			21017: outdata = 32'd44519;
			21018: outdata = 32'd44518;
			21019: outdata = 32'd44517;
			21020: outdata = 32'd44516;
			21021: outdata = 32'd44515;
			21022: outdata = 32'd44514;
			21023: outdata = 32'd44513;
			21024: outdata = 32'd44512;
			21025: outdata = 32'd44511;
			21026: outdata = 32'd44510;
			21027: outdata = 32'd44509;
			21028: outdata = 32'd44508;
			21029: outdata = 32'd44507;
			21030: outdata = 32'd44506;
			21031: outdata = 32'd44505;
			21032: outdata = 32'd44504;
			21033: outdata = 32'd44503;
			21034: outdata = 32'd44502;
			21035: outdata = 32'd44501;
			21036: outdata = 32'd44500;
			21037: outdata = 32'd44499;
			21038: outdata = 32'd44498;
			21039: outdata = 32'd44497;
			21040: outdata = 32'd44496;
			21041: outdata = 32'd44495;
			21042: outdata = 32'd44494;
			21043: outdata = 32'd44493;
			21044: outdata = 32'd44492;
			21045: outdata = 32'd44491;
			21046: outdata = 32'd44490;
			21047: outdata = 32'd44489;
			21048: outdata = 32'd44488;
			21049: outdata = 32'd44487;
			21050: outdata = 32'd44486;
			21051: outdata = 32'd44485;
			21052: outdata = 32'd44484;
			21053: outdata = 32'd44483;
			21054: outdata = 32'd44482;
			21055: outdata = 32'd44481;
			21056: outdata = 32'd44480;
			21057: outdata = 32'd44479;
			21058: outdata = 32'd44478;
			21059: outdata = 32'd44477;
			21060: outdata = 32'd44476;
			21061: outdata = 32'd44475;
			21062: outdata = 32'd44474;
			21063: outdata = 32'd44473;
			21064: outdata = 32'd44472;
			21065: outdata = 32'd44471;
			21066: outdata = 32'd44470;
			21067: outdata = 32'd44469;
			21068: outdata = 32'd44468;
			21069: outdata = 32'd44467;
			21070: outdata = 32'd44466;
			21071: outdata = 32'd44465;
			21072: outdata = 32'd44464;
			21073: outdata = 32'd44463;
			21074: outdata = 32'd44462;
			21075: outdata = 32'd44461;
			21076: outdata = 32'd44460;
			21077: outdata = 32'd44459;
			21078: outdata = 32'd44458;
			21079: outdata = 32'd44457;
			21080: outdata = 32'd44456;
			21081: outdata = 32'd44455;
			21082: outdata = 32'd44454;
			21083: outdata = 32'd44453;
			21084: outdata = 32'd44452;
			21085: outdata = 32'd44451;
			21086: outdata = 32'd44450;
			21087: outdata = 32'd44449;
			21088: outdata = 32'd44448;
			21089: outdata = 32'd44447;
			21090: outdata = 32'd44446;
			21091: outdata = 32'd44445;
			21092: outdata = 32'd44444;
			21093: outdata = 32'd44443;
			21094: outdata = 32'd44442;
			21095: outdata = 32'd44441;
			21096: outdata = 32'd44440;
			21097: outdata = 32'd44439;
			21098: outdata = 32'd44438;
			21099: outdata = 32'd44437;
			21100: outdata = 32'd44436;
			21101: outdata = 32'd44435;
			21102: outdata = 32'd44434;
			21103: outdata = 32'd44433;
			21104: outdata = 32'd44432;
			21105: outdata = 32'd44431;
			21106: outdata = 32'd44430;
			21107: outdata = 32'd44429;
			21108: outdata = 32'd44428;
			21109: outdata = 32'd44427;
			21110: outdata = 32'd44426;
			21111: outdata = 32'd44425;
			21112: outdata = 32'd44424;
			21113: outdata = 32'd44423;
			21114: outdata = 32'd44422;
			21115: outdata = 32'd44421;
			21116: outdata = 32'd44420;
			21117: outdata = 32'd44419;
			21118: outdata = 32'd44418;
			21119: outdata = 32'd44417;
			21120: outdata = 32'd44416;
			21121: outdata = 32'd44415;
			21122: outdata = 32'd44414;
			21123: outdata = 32'd44413;
			21124: outdata = 32'd44412;
			21125: outdata = 32'd44411;
			21126: outdata = 32'd44410;
			21127: outdata = 32'd44409;
			21128: outdata = 32'd44408;
			21129: outdata = 32'd44407;
			21130: outdata = 32'd44406;
			21131: outdata = 32'd44405;
			21132: outdata = 32'd44404;
			21133: outdata = 32'd44403;
			21134: outdata = 32'd44402;
			21135: outdata = 32'd44401;
			21136: outdata = 32'd44400;
			21137: outdata = 32'd44399;
			21138: outdata = 32'd44398;
			21139: outdata = 32'd44397;
			21140: outdata = 32'd44396;
			21141: outdata = 32'd44395;
			21142: outdata = 32'd44394;
			21143: outdata = 32'd44393;
			21144: outdata = 32'd44392;
			21145: outdata = 32'd44391;
			21146: outdata = 32'd44390;
			21147: outdata = 32'd44389;
			21148: outdata = 32'd44388;
			21149: outdata = 32'd44387;
			21150: outdata = 32'd44386;
			21151: outdata = 32'd44385;
			21152: outdata = 32'd44384;
			21153: outdata = 32'd44383;
			21154: outdata = 32'd44382;
			21155: outdata = 32'd44381;
			21156: outdata = 32'd44380;
			21157: outdata = 32'd44379;
			21158: outdata = 32'd44378;
			21159: outdata = 32'd44377;
			21160: outdata = 32'd44376;
			21161: outdata = 32'd44375;
			21162: outdata = 32'd44374;
			21163: outdata = 32'd44373;
			21164: outdata = 32'd44372;
			21165: outdata = 32'd44371;
			21166: outdata = 32'd44370;
			21167: outdata = 32'd44369;
			21168: outdata = 32'd44368;
			21169: outdata = 32'd44367;
			21170: outdata = 32'd44366;
			21171: outdata = 32'd44365;
			21172: outdata = 32'd44364;
			21173: outdata = 32'd44363;
			21174: outdata = 32'd44362;
			21175: outdata = 32'd44361;
			21176: outdata = 32'd44360;
			21177: outdata = 32'd44359;
			21178: outdata = 32'd44358;
			21179: outdata = 32'd44357;
			21180: outdata = 32'd44356;
			21181: outdata = 32'd44355;
			21182: outdata = 32'd44354;
			21183: outdata = 32'd44353;
			21184: outdata = 32'd44352;
			21185: outdata = 32'd44351;
			21186: outdata = 32'd44350;
			21187: outdata = 32'd44349;
			21188: outdata = 32'd44348;
			21189: outdata = 32'd44347;
			21190: outdata = 32'd44346;
			21191: outdata = 32'd44345;
			21192: outdata = 32'd44344;
			21193: outdata = 32'd44343;
			21194: outdata = 32'd44342;
			21195: outdata = 32'd44341;
			21196: outdata = 32'd44340;
			21197: outdata = 32'd44339;
			21198: outdata = 32'd44338;
			21199: outdata = 32'd44337;
			21200: outdata = 32'd44336;
			21201: outdata = 32'd44335;
			21202: outdata = 32'd44334;
			21203: outdata = 32'd44333;
			21204: outdata = 32'd44332;
			21205: outdata = 32'd44331;
			21206: outdata = 32'd44330;
			21207: outdata = 32'd44329;
			21208: outdata = 32'd44328;
			21209: outdata = 32'd44327;
			21210: outdata = 32'd44326;
			21211: outdata = 32'd44325;
			21212: outdata = 32'd44324;
			21213: outdata = 32'd44323;
			21214: outdata = 32'd44322;
			21215: outdata = 32'd44321;
			21216: outdata = 32'd44320;
			21217: outdata = 32'd44319;
			21218: outdata = 32'd44318;
			21219: outdata = 32'd44317;
			21220: outdata = 32'd44316;
			21221: outdata = 32'd44315;
			21222: outdata = 32'd44314;
			21223: outdata = 32'd44313;
			21224: outdata = 32'd44312;
			21225: outdata = 32'd44311;
			21226: outdata = 32'd44310;
			21227: outdata = 32'd44309;
			21228: outdata = 32'd44308;
			21229: outdata = 32'd44307;
			21230: outdata = 32'd44306;
			21231: outdata = 32'd44305;
			21232: outdata = 32'd44304;
			21233: outdata = 32'd44303;
			21234: outdata = 32'd44302;
			21235: outdata = 32'd44301;
			21236: outdata = 32'd44300;
			21237: outdata = 32'd44299;
			21238: outdata = 32'd44298;
			21239: outdata = 32'd44297;
			21240: outdata = 32'd44296;
			21241: outdata = 32'd44295;
			21242: outdata = 32'd44294;
			21243: outdata = 32'd44293;
			21244: outdata = 32'd44292;
			21245: outdata = 32'd44291;
			21246: outdata = 32'd44290;
			21247: outdata = 32'd44289;
			21248: outdata = 32'd44288;
			21249: outdata = 32'd44287;
			21250: outdata = 32'd44286;
			21251: outdata = 32'd44285;
			21252: outdata = 32'd44284;
			21253: outdata = 32'd44283;
			21254: outdata = 32'd44282;
			21255: outdata = 32'd44281;
			21256: outdata = 32'd44280;
			21257: outdata = 32'd44279;
			21258: outdata = 32'd44278;
			21259: outdata = 32'd44277;
			21260: outdata = 32'd44276;
			21261: outdata = 32'd44275;
			21262: outdata = 32'd44274;
			21263: outdata = 32'd44273;
			21264: outdata = 32'd44272;
			21265: outdata = 32'd44271;
			21266: outdata = 32'd44270;
			21267: outdata = 32'd44269;
			21268: outdata = 32'd44268;
			21269: outdata = 32'd44267;
			21270: outdata = 32'd44266;
			21271: outdata = 32'd44265;
			21272: outdata = 32'd44264;
			21273: outdata = 32'd44263;
			21274: outdata = 32'd44262;
			21275: outdata = 32'd44261;
			21276: outdata = 32'd44260;
			21277: outdata = 32'd44259;
			21278: outdata = 32'd44258;
			21279: outdata = 32'd44257;
			21280: outdata = 32'd44256;
			21281: outdata = 32'd44255;
			21282: outdata = 32'd44254;
			21283: outdata = 32'd44253;
			21284: outdata = 32'd44252;
			21285: outdata = 32'd44251;
			21286: outdata = 32'd44250;
			21287: outdata = 32'd44249;
			21288: outdata = 32'd44248;
			21289: outdata = 32'd44247;
			21290: outdata = 32'd44246;
			21291: outdata = 32'd44245;
			21292: outdata = 32'd44244;
			21293: outdata = 32'd44243;
			21294: outdata = 32'd44242;
			21295: outdata = 32'd44241;
			21296: outdata = 32'd44240;
			21297: outdata = 32'd44239;
			21298: outdata = 32'd44238;
			21299: outdata = 32'd44237;
			21300: outdata = 32'd44236;
			21301: outdata = 32'd44235;
			21302: outdata = 32'd44234;
			21303: outdata = 32'd44233;
			21304: outdata = 32'd44232;
			21305: outdata = 32'd44231;
			21306: outdata = 32'd44230;
			21307: outdata = 32'd44229;
			21308: outdata = 32'd44228;
			21309: outdata = 32'd44227;
			21310: outdata = 32'd44226;
			21311: outdata = 32'd44225;
			21312: outdata = 32'd44224;
			21313: outdata = 32'd44223;
			21314: outdata = 32'd44222;
			21315: outdata = 32'd44221;
			21316: outdata = 32'd44220;
			21317: outdata = 32'd44219;
			21318: outdata = 32'd44218;
			21319: outdata = 32'd44217;
			21320: outdata = 32'd44216;
			21321: outdata = 32'd44215;
			21322: outdata = 32'd44214;
			21323: outdata = 32'd44213;
			21324: outdata = 32'd44212;
			21325: outdata = 32'd44211;
			21326: outdata = 32'd44210;
			21327: outdata = 32'd44209;
			21328: outdata = 32'd44208;
			21329: outdata = 32'd44207;
			21330: outdata = 32'd44206;
			21331: outdata = 32'd44205;
			21332: outdata = 32'd44204;
			21333: outdata = 32'd44203;
			21334: outdata = 32'd44202;
			21335: outdata = 32'd44201;
			21336: outdata = 32'd44200;
			21337: outdata = 32'd44199;
			21338: outdata = 32'd44198;
			21339: outdata = 32'd44197;
			21340: outdata = 32'd44196;
			21341: outdata = 32'd44195;
			21342: outdata = 32'd44194;
			21343: outdata = 32'd44193;
			21344: outdata = 32'd44192;
			21345: outdata = 32'd44191;
			21346: outdata = 32'd44190;
			21347: outdata = 32'd44189;
			21348: outdata = 32'd44188;
			21349: outdata = 32'd44187;
			21350: outdata = 32'd44186;
			21351: outdata = 32'd44185;
			21352: outdata = 32'd44184;
			21353: outdata = 32'd44183;
			21354: outdata = 32'd44182;
			21355: outdata = 32'd44181;
			21356: outdata = 32'd44180;
			21357: outdata = 32'd44179;
			21358: outdata = 32'd44178;
			21359: outdata = 32'd44177;
			21360: outdata = 32'd44176;
			21361: outdata = 32'd44175;
			21362: outdata = 32'd44174;
			21363: outdata = 32'd44173;
			21364: outdata = 32'd44172;
			21365: outdata = 32'd44171;
			21366: outdata = 32'd44170;
			21367: outdata = 32'd44169;
			21368: outdata = 32'd44168;
			21369: outdata = 32'd44167;
			21370: outdata = 32'd44166;
			21371: outdata = 32'd44165;
			21372: outdata = 32'd44164;
			21373: outdata = 32'd44163;
			21374: outdata = 32'd44162;
			21375: outdata = 32'd44161;
			21376: outdata = 32'd44160;
			21377: outdata = 32'd44159;
			21378: outdata = 32'd44158;
			21379: outdata = 32'd44157;
			21380: outdata = 32'd44156;
			21381: outdata = 32'd44155;
			21382: outdata = 32'd44154;
			21383: outdata = 32'd44153;
			21384: outdata = 32'd44152;
			21385: outdata = 32'd44151;
			21386: outdata = 32'd44150;
			21387: outdata = 32'd44149;
			21388: outdata = 32'd44148;
			21389: outdata = 32'd44147;
			21390: outdata = 32'd44146;
			21391: outdata = 32'd44145;
			21392: outdata = 32'd44144;
			21393: outdata = 32'd44143;
			21394: outdata = 32'd44142;
			21395: outdata = 32'd44141;
			21396: outdata = 32'd44140;
			21397: outdata = 32'd44139;
			21398: outdata = 32'd44138;
			21399: outdata = 32'd44137;
			21400: outdata = 32'd44136;
			21401: outdata = 32'd44135;
			21402: outdata = 32'd44134;
			21403: outdata = 32'd44133;
			21404: outdata = 32'd44132;
			21405: outdata = 32'd44131;
			21406: outdata = 32'd44130;
			21407: outdata = 32'd44129;
			21408: outdata = 32'd44128;
			21409: outdata = 32'd44127;
			21410: outdata = 32'd44126;
			21411: outdata = 32'd44125;
			21412: outdata = 32'd44124;
			21413: outdata = 32'd44123;
			21414: outdata = 32'd44122;
			21415: outdata = 32'd44121;
			21416: outdata = 32'd44120;
			21417: outdata = 32'd44119;
			21418: outdata = 32'd44118;
			21419: outdata = 32'd44117;
			21420: outdata = 32'd44116;
			21421: outdata = 32'd44115;
			21422: outdata = 32'd44114;
			21423: outdata = 32'd44113;
			21424: outdata = 32'd44112;
			21425: outdata = 32'd44111;
			21426: outdata = 32'd44110;
			21427: outdata = 32'd44109;
			21428: outdata = 32'd44108;
			21429: outdata = 32'd44107;
			21430: outdata = 32'd44106;
			21431: outdata = 32'd44105;
			21432: outdata = 32'd44104;
			21433: outdata = 32'd44103;
			21434: outdata = 32'd44102;
			21435: outdata = 32'd44101;
			21436: outdata = 32'd44100;
			21437: outdata = 32'd44099;
			21438: outdata = 32'd44098;
			21439: outdata = 32'd44097;
			21440: outdata = 32'd44096;
			21441: outdata = 32'd44095;
			21442: outdata = 32'd44094;
			21443: outdata = 32'd44093;
			21444: outdata = 32'd44092;
			21445: outdata = 32'd44091;
			21446: outdata = 32'd44090;
			21447: outdata = 32'd44089;
			21448: outdata = 32'd44088;
			21449: outdata = 32'd44087;
			21450: outdata = 32'd44086;
			21451: outdata = 32'd44085;
			21452: outdata = 32'd44084;
			21453: outdata = 32'd44083;
			21454: outdata = 32'd44082;
			21455: outdata = 32'd44081;
			21456: outdata = 32'd44080;
			21457: outdata = 32'd44079;
			21458: outdata = 32'd44078;
			21459: outdata = 32'd44077;
			21460: outdata = 32'd44076;
			21461: outdata = 32'd44075;
			21462: outdata = 32'd44074;
			21463: outdata = 32'd44073;
			21464: outdata = 32'd44072;
			21465: outdata = 32'd44071;
			21466: outdata = 32'd44070;
			21467: outdata = 32'd44069;
			21468: outdata = 32'd44068;
			21469: outdata = 32'd44067;
			21470: outdata = 32'd44066;
			21471: outdata = 32'd44065;
			21472: outdata = 32'd44064;
			21473: outdata = 32'd44063;
			21474: outdata = 32'd44062;
			21475: outdata = 32'd44061;
			21476: outdata = 32'd44060;
			21477: outdata = 32'd44059;
			21478: outdata = 32'd44058;
			21479: outdata = 32'd44057;
			21480: outdata = 32'd44056;
			21481: outdata = 32'd44055;
			21482: outdata = 32'd44054;
			21483: outdata = 32'd44053;
			21484: outdata = 32'd44052;
			21485: outdata = 32'd44051;
			21486: outdata = 32'd44050;
			21487: outdata = 32'd44049;
			21488: outdata = 32'd44048;
			21489: outdata = 32'd44047;
			21490: outdata = 32'd44046;
			21491: outdata = 32'd44045;
			21492: outdata = 32'd44044;
			21493: outdata = 32'd44043;
			21494: outdata = 32'd44042;
			21495: outdata = 32'd44041;
			21496: outdata = 32'd44040;
			21497: outdata = 32'd44039;
			21498: outdata = 32'd44038;
			21499: outdata = 32'd44037;
			21500: outdata = 32'd44036;
			21501: outdata = 32'd44035;
			21502: outdata = 32'd44034;
			21503: outdata = 32'd44033;
			21504: outdata = 32'd44032;
			21505: outdata = 32'd44031;
			21506: outdata = 32'd44030;
			21507: outdata = 32'd44029;
			21508: outdata = 32'd44028;
			21509: outdata = 32'd44027;
			21510: outdata = 32'd44026;
			21511: outdata = 32'd44025;
			21512: outdata = 32'd44024;
			21513: outdata = 32'd44023;
			21514: outdata = 32'd44022;
			21515: outdata = 32'd44021;
			21516: outdata = 32'd44020;
			21517: outdata = 32'd44019;
			21518: outdata = 32'd44018;
			21519: outdata = 32'd44017;
			21520: outdata = 32'd44016;
			21521: outdata = 32'd44015;
			21522: outdata = 32'd44014;
			21523: outdata = 32'd44013;
			21524: outdata = 32'd44012;
			21525: outdata = 32'd44011;
			21526: outdata = 32'd44010;
			21527: outdata = 32'd44009;
			21528: outdata = 32'd44008;
			21529: outdata = 32'd44007;
			21530: outdata = 32'd44006;
			21531: outdata = 32'd44005;
			21532: outdata = 32'd44004;
			21533: outdata = 32'd44003;
			21534: outdata = 32'd44002;
			21535: outdata = 32'd44001;
			21536: outdata = 32'd44000;
			21537: outdata = 32'd43999;
			21538: outdata = 32'd43998;
			21539: outdata = 32'd43997;
			21540: outdata = 32'd43996;
			21541: outdata = 32'd43995;
			21542: outdata = 32'd43994;
			21543: outdata = 32'd43993;
			21544: outdata = 32'd43992;
			21545: outdata = 32'd43991;
			21546: outdata = 32'd43990;
			21547: outdata = 32'd43989;
			21548: outdata = 32'd43988;
			21549: outdata = 32'd43987;
			21550: outdata = 32'd43986;
			21551: outdata = 32'd43985;
			21552: outdata = 32'd43984;
			21553: outdata = 32'd43983;
			21554: outdata = 32'd43982;
			21555: outdata = 32'd43981;
			21556: outdata = 32'd43980;
			21557: outdata = 32'd43979;
			21558: outdata = 32'd43978;
			21559: outdata = 32'd43977;
			21560: outdata = 32'd43976;
			21561: outdata = 32'd43975;
			21562: outdata = 32'd43974;
			21563: outdata = 32'd43973;
			21564: outdata = 32'd43972;
			21565: outdata = 32'd43971;
			21566: outdata = 32'd43970;
			21567: outdata = 32'd43969;
			21568: outdata = 32'd43968;
			21569: outdata = 32'd43967;
			21570: outdata = 32'd43966;
			21571: outdata = 32'd43965;
			21572: outdata = 32'd43964;
			21573: outdata = 32'd43963;
			21574: outdata = 32'd43962;
			21575: outdata = 32'd43961;
			21576: outdata = 32'd43960;
			21577: outdata = 32'd43959;
			21578: outdata = 32'd43958;
			21579: outdata = 32'd43957;
			21580: outdata = 32'd43956;
			21581: outdata = 32'd43955;
			21582: outdata = 32'd43954;
			21583: outdata = 32'd43953;
			21584: outdata = 32'd43952;
			21585: outdata = 32'd43951;
			21586: outdata = 32'd43950;
			21587: outdata = 32'd43949;
			21588: outdata = 32'd43948;
			21589: outdata = 32'd43947;
			21590: outdata = 32'd43946;
			21591: outdata = 32'd43945;
			21592: outdata = 32'd43944;
			21593: outdata = 32'd43943;
			21594: outdata = 32'd43942;
			21595: outdata = 32'd43941;
			21596: outdata = 32'd43940;
			21597: outdata = 32'd43939;
			21598: outdata = 32'd43938;
			21599: outdata = 32'd43937;
			21600: outdata = 32'd43936;
			21601: outdata = 32'd43935;
			21602: outdata = 32'd43934;
			21603: outdata = 32'd43933;
			21604: outdata = 32'd43932;
			21605: outdata = 32'd43931;
			21606: outdata = 32'd43930;
			21607: outdata = 32'd43929;
			21608: outdata = 32'd43928;
			21609: outdata = 32'd43927;
			21610: outdata = 32'd43926;
			21611: outdata = 32'd43925;
			21612: outdata = 32'd43924;
			21613: outdata = 32'd43923;
			21614: outdata = 32'd43922;
			21615: outdata = 32'd43921;
			21616: outdata = 32'd43920;
			21617: outdata = 32'd43919;
			21618: outdata = 32'd43918;
			21619: outdata = 32'd43917;
			21620: outdata = 32'd43916;
			21621: outdata = 32'd43915;
			21622: outdata = 32'd43914;
			21623: outdata = 32'd43913;
			21624: outdata = 32'd43912;
			21625: outdata = 32'd43911;
			21626: outdata = 32'd43910;
			21627: outdata = 32'd43909;
			21628: outdata = 32'd43908;
			21629: outdata = 32'd43907;
			21630: outdata = 32'd43906;
			21631: outdata = 32'd43905;
			21632: outdata = 32'd43904;
			21633: outdata = 32'd43903;
			21634: outdata = 32'd43902;
			21635: outdata = 32'd43901;
			21636: outdata = 32'd43900;
			21637: outdata = 32'd43899;
			21638: outdata = 32'd43898;
			21639: outdata = 32'd43897;
			21640: outdata = 32'd43896;
			21641: outdata = 32'd43895;
			21642: outdata = 32'd43894;
			21643: outdata = 32'd43893;
			21644: outdata = 32'd43892;
			21645: outdata = 32'd43891;
			21646: outdata = 32'd43890;
			21647: outdata = 32'd43889;
			21648: outdata = 32'd43888;
			21649: outdata = 32'd43887;
			21650: outdata = 32'd43886;
			21651: outdata = 32'd43885;
			21652: outdata = 32'd43884;
			21653: outdata = 32'd43883;
			21654: outdata = 32'd43882;
			21655: outdata = 32'd43881;
			21656: outdata = 32'd43880;
			21657: outdata = 32'd43879;
			21658: outdata = 32'd43878;
			21659: outdata = 32'd43877;
			21660: outdata = 32'd43876;
			21661: outdata = 32'd43875;
			21662: outdata = 32'd43874;
			21663: outdata = 32'd43873;
			21664: outdata = 32'd43872;
			21665: outdata = 32'd43871;
			21666: outdata = 32'd43870;
			21667: outdata = 32'd43869;
			21668: outdata = 32'd43868;
			21669: outdata = 32'd43867;
			21670: outdata = 32'd43866;
			21671: outdata = 32'd43865;
			21672: outdata = 32'd43864;
			21673: outdata = 32'd43863;
			21674: outdata = 32'd43862;
			21675: outdata = 32'd43861;
			21676: outdata = 32'd43860;
			21677: outdata = 32'd43859;
			21678: outdata = 32'd43858;
			21679: outdata = 32'd43857;
			21680: outdata = 32'd43856;
			21681: outdata = 32'd43855;
			21682: outdata = 32'd43854;
			21683: outdata = 32'd43853;
			21684: outdata = 32'd43852;
			21685: outdata = 32'd43851;
			21686: outdata = 32'd43850;
			21687: outdata = 32'd43849;
			21688: outdata = 32'd43848;
			21689: outdata = 32'd43847;
			21690: outdata = 32'd43846;
			21691: outdata = 32'd43845;
			21692: outdata = 32'd43844;
			21693: outdata = 32'd43843;
			21694: outdata = 32'd43842;
			21695: outdata = 32'd43841;
			21696: outdata = 32'd43840;
			21697: outdata = 32'd43839;
			21698: outdata = 32'd43838;
			21699: outdata = 32'd43837;
			21700: outdata = 32'd43836;
			21701: outdata = 32'd43835;
			21702: outdata = 32'd43834;
			21703: outdata = 32'd43833;
			21704: outdata = 32'd43832;
			21705: outdata = 32'd43831;
			21706: outdata = 32'd43830;
			21707: outdata = 32'd43829;
			21708: outdata = 32'd43828;
			21709: outdata = 32'd43827;
			21710: outdata = 32'd43826;
			21711: outdata = 32'd43825;
			21712: outdata = 32'd43824;
			21713: outdata = 32'd43823;
			21714: outdata = 32'd43822;
			21715: outdata = 32'd43821;
			21716: outdata = 32'd43820;
			21717: outdata = 32'd43819;
			21718: outdata = 32'd43818;
			21719: outdata = 32'd43817;
			21720: outdata = 32'd43816;
			21721: outdata = 32'd43815;
			21722: outdata = 32'd43814;
			21723: outdata = 32'd43813;
			21724: outdata = 32'd43812;
			21725: outdata = 32'd43811;
			21726: outdata = 32'd43810;
			21727: outdata = 32'd43809;
			21728: outdata = 32'd43808;
			21729: outdata = 32'd43807;
			21730: outdata = 32'd43806;
			21731: outdata = 32'd43805;
			21732: outdata = 32'd43804;
			21733: outdata = 32'd43803;
			21734: outdata = 32'd43802;
			21735: outdata = 32'd43801;
			21736: outdata = 32'd43800;
			21737: outdata = 32'd43799;
			21738: outdata = 32'd43798;
			21739: outdata = 32'd43797;
			21740: outdata = 32'd43796;
			21741: outdata = 32'd43795;
			21742: outdata = 32'd43794;
			21743: outdata = 32'd43793;
			21744: outdata = 32'd43792;
			21745: outdata = 32'd43791;
			21746: outdata = 32'd43790;
			21747: outdata = 32'd43789;
			21748: outdata = 32'd43788;
			21749: outdata = 32'd43787;
			21750: outdata = 32'd43786;
			21751: outdata = 32'd43785;
			21752: outdata = 32'd43784;
			21753: outdata = 32'd43783;
			21754: outdata = 32'd43782;
			21755: outdata = 32'd43781;
			21756: outdata = 32'd43780;
			21757: outdata = 32'd43779;
			21758: outdata = 32'd43778;
			21759: outdata = 32'd43777;
			21760: outdata = 32'd43776;
			21761: outdata = 32'd43775;
			21762: outdata = 32'd43774;
			21763: outdata = 32'd43773;
			21764: outdata = 32'd43772;
			21765: outdata = 32'd43771;
			21766: outdata = 32'd43770;
			21767: outdata = 32'd43769;
			21768: outdata = 32'd43768;
			21769: outdata = 32'd43767;
			21770: outdata = 32'd43766;
			21771: outdata = 32'd43765;
			21772: outdata = 32'd43764;
			21773: outdata = 32'd43763;
			21774: outdata = 32'd43762;
			21775: outdata = 32'd43761;
			21776: outdata = 32'd43760;
			21777: outdata = 32'd43759;
			21778: outdata = 32'd43758;
			21779: outdata = 32'd43757;
			21780: outdata = 32'd43756;
			21781: outdata = 32'd43755;
			21782: outdata = 32'd43754;
			21783: outdata = 32'd43753;
			21784: outdata = 32'd43752;
			21785: outdata = 32'd43751;
			21786: outdata = 32'd43750;
			21787: outdata = 32'd43749;
			21788: outdata = 32'd43748;
			21789: outdata = 32'd43747;
			21790: outdata = 32'd43746;
			21791: outdata = 32'd43745;
			21792: outdata = 32'd43744;
			21793: outdata = 32'd43743;
			21794: outdata = 32'd43742;
			21795: outdata = 32'd43741;
			21796: outdata = 32'd43740;
			21797: outdata = 32'd43739;
			21798: outdata = 32'd43738;
			21799: outdata = 32'd43737;
			21800: outdata = 32'd43736;
			21801: outdata = 32'd43735;
			21802: outdata = 32'd43734;
			21803: outdata = 32'd43733;
			21804: outdata = 32'd43732;
			21805: outdata = 32'd43731;
			21806: outdata = 32'd43730;
			21807: outdata = 32'd43729;
			21808: outdata = 32'd43728;
			21809: outdata = 32'd43727;
			21810: outdata = 32'd43726;
			21811: outdata = 32'd43725;
			21812: outdata = 32'd43724;
			21813: outdata = 32'd43723;
			21814: outdata = 32'd43722;
			21815: outdata = 32'd43721;
			21816: outdata = 32'd43720;
			21817: outdata = 32'd43719;
			21818: outdata = 32'd43718;
			21819: outdata = 32'd43717;
			21820: outdata = 32'd43716;
			21821: outdata = 32'd43715;
			21822: outdata = 32'd43714;
			21823: outdata = 32'd43713;
			21824: outdata = 32'd43712;
			21825: outdata = 32'd43711;
			21826: outdata = 32'd43710;
			21827: outdata = 32'd43709;
			21828: outdata = 32'd43708;
			21829: outdata = 32'd43707;
			21830: outdata = 32'd43706;
			21831: outdata = 32'd43705;
			21832: outdata = 32'd43704;
			21833: outdata = 32'd43703;
			21834: outdata = 32'd43702;
			21835: outdata = 32'd43701;
			21836: outdata = 32'd43700;
			21837: outdata = 32'd43699;
			21838: outdata = 32'd43698;
			21839: outdata = 32'd43697;
			21840: outdata = 32'd43696;
			21841: outdata = 32'd43695;
			21842: outdata = 32'd43694;
			21843: outdata = 32'd43693;
			21844: outdata = 32'd43692;
			21845: outdata = 32'd43691;
			21846: outdata = 32'd43690;
			21847: outdata = 32'd43689;
			21848: outdata = 32'd43688;
			21849: outdata = 32'd43687;
			21850: outdata = 32'd43686;
			21851: outdata = 32'd43685;
			21852: outdata = 32'd43684;
			21853: outdata = 32'd43683;
			21854: outdata = 32'd43682;
			21855: outdata = 32'd43681;
			21856: outdata = 32'd43680;
			21857: outdata = 32'd43679;
			21858: outdata = 32'd43678;
			21859: outdata = 32'd43677;
			21860: outdata = 32'd43676;
			21861: outdata = 32'd43675;
			21862: outdata = 32'd43674;
			21863: outdata = 32'd43673;
			21864: outdata = 32'd43672;
			21865: outdata = 32'd43671;
			21866: outdata = 32'd43670;
			21867: outdata = 32'd43669;
			21868: outdata = 32'd43668;
			21869: outdata = 32'd43667;
			21870: outdata = 32'd43666;
			21871: outdata = 32'd43665;
			21872: outdata = 32'd43664;
			21873: outdata = 32'd43663;
			21874: outdata = 32'd43662;
			21875: outdata = 32'd43661;
			21876: outdata = 32'd43660;
			21877: outdata = 32'd43659;
			21878: outdata = 32'd43658;
			21879: outdata = 32'd43657;
			21880: outdata = 32'd43656;
			21881: outdata = 32'd43655;
			21882: outdata = 32'd43654;
			21883: outdata = 32'd43653;
			21884: outdata = 32'd43652;
			21885: outdata = 32'd43651;
			21886: outdata = 32'd43650;
			21887: outdata = 32'd43649;
			21888: outdata = 32'd43648;
			21889: outdata = 32'd43647;
			21890: outdata = 32'd43646;
			21891: outdata = 32'd43645;
			21892: outdata = 32'd43644;
			21893: outdata = 32'd43643;
			21894: outdata = 32'd43642;
			21895: outdata = 32'd43641;
			21896: outdata = 32'd43640;
			21897: outdata = 32'd43639;
			21898: outdata = 32'd43638;
			21899: outdata = 32'd43637;
			21900: outdata = 32'd43636;
			21901: outdata = 32'd43635;
			21902: outdata = 32'd43634;
			21903: outdata = 32'd43633;
			21904: outdata = 32'd43632;
			21905: outdata = 32'd43631;
			21906: outdata = 32'd43630;
			21907: outdata = 32'd43629;
			21908: outdata = 32'd43628;
			21909: outdata = 32'd43627;
			21910: outdata = 32'd43626;
			21911: outdata = 32'd43625;
			21912: outdata = 32'd43624;
			21913: outdata = 32'd43623;
			21914: outdata = 32'd43622;
			21915: outdata = 32'd43621;
			21916: outdata = 32'd43620;
			21917: outdata = 32'd43619;
			21918: outdata = 32'd43618;
			21919: outdata = 32'd43617;
			21920: outdata = 32'd43616;
			21921: outdata = 32'd43615;
			21922: outdata = 32'd43614;
			21923: outdata = 32'd43613;
			21924: outdata = 32'd43612;
			21925: outdata = 32'd43611;
			21926: outdata = 32'd43610;
			21927: outdata = 32'd43609;
			21928: outdata = 32'd43608;
			21929: outdata = 32'd43607;
			21930: outdata = 32'd43606;
			21931: outdata = 32'd43605;
			21932: outdata = 32'd43604;
			21933: outdata = 32'd43603;
			21934: outdata = 32'd43602;
			21935: outdata = 32'd43601;
			21936: outdata = 32'd43600;
			21937: outdata = 32'd43599;
			21938: outdata = 32'd43598;
			21939: outdata = 32'd43597;
			21940: outdata = 32'd43596;
			21941: outdata = 32'd43595;
			21942: outdata = 32'd43594;
			21943: outdata = 32'd43593;
			21944: outdata = 32'd43592;
			21945: outdata = 32'd43591;
			21946: outdata = 32'd43590;
			21947: outdata = 32'd43589;
			21948: outdata = 32'd43588;
			21949: outdata = 32'd43587;
			21950: outdata = 32'd43586;
			21951: outdata = 32'd43585;
			21952: outdata = 32'd43584;
			21953: outdata = 32'd43583;
			21954: outdata = 32'd43582;
			21955: outdata = 32'd43581;
			21956: outdata = 32'd43580;
			21957: outdata = 32'd43579;
			21958: outdata = 32'd43578;
			21959: outdata = 32'd43577;
			21960: outdata = 32'd43576;
			21961: outdata = 32'd43575;
			21962: outdata = 32'd43574;
			21963: outdata = 32'd43573;
			21964: outdata = 32'd43572;
			21965: outdata = 32'd43571;
			21966: outdata = 32'd43570;
			21967: outdata = 32'd43569;
			21968: outdata = 32'd43568;
			21969: outdata = 32'd43567;
			21970: outdata = 32'd43566;
			21971: outdata = 32'd43565;
			21972: outdata = 32'd43564;
			21973: outdata = 32'd43563;
			21974: outdata = 32'd43562;
			21975: outdata = 32'd43561;
			21976: outdata = 32'd43560;
			21977: outdata = 32'd43559;
			21978: outdata = 32'd43558;
			21979: outdata = 32'd43557;
			21980: outdata = 32'd43556;
			21981: outdata = 32'd43555;
			21982: outdata = 32'd43554;
			21983: outdata = 32'd43553;
			21984: outdata = 32'd43552;
			21985: outdata = 32'd43551;
			21986: outdata = 32'd43550;
			21987: outdata = 32'd43549;
			21988: outdata = 32'd43548;
			21989: outdata = 32'd43547;
			21990: outdata = 32'd43546;
			21991: outdata = 32'd43545;
			21992: outdata = 32'd43544;
			21993: outdata = 32'd43543;
			21994: outdata = 32'd43542;
			21995: outdata = 32'd43541;
			21996: outdata = 32'd43540;
			21997: outdata = 32'd43539;
			21998: outdata = 32'd43538;
			21999: outdata = 32'd43537;
			22000: outdata = 32'd43536;
			22001: outdata = 32'd43535;
			22002: outdata = 32'd43534;
			22003: outdata = 32'd43533;
			22004: outdata = 32'd43532;
			22005: outdata = 32'd43531;
			22006: outdata = 32'd43530;
			22007: outdata = 32'd43529;
			22008: outdata = 32'd43528;
			22009: outdata = 32'd43527;
			22010: outdata = 32'd43526;
			22011: outdata = 32'd43525;
			22012: outdata = 32'd43524;
			22013: outdata = 32'd43523;
			22014: outdata = 32'd43522;
			22015: outdata = 32'd43521;
			22016: outdata = 32'd43520;
			22017: outdata = 32'd43519;
			22018: outdata = 32'd43518;
			22019: outdata = 32'd43517;
			22020: outdata = 32'd43516;
			22021: outdata = 32'd43515;
			22022: outdata = 32'd43514;
			22023: outdata = 32'd43513;
			22024: outdata = 32'd43512;
			22025: outdata = 32'd43511;
			22026: outdata = 32'd43510;
			22027: outdata = 32'd43509;
			22028: outdata = 32'd43508;
			22029: outdata = 32'd43507;
			22030: outdata = 32'd43506;
			22031: outdata = 32'd43505;
			22032: outdata = 32'd43504;
			22033: outdata = 32'd43503;
			22034: outdata = 32'd43502;
			22035: outdata = 32'd43501;
			22036: outdata = 32'd43500;
			22037: outdata = 32'd43499;
			22038: outdata = 32'd43498;
			22039: outdata = 32'd43497;
			22040: outdata = 32'd43496;
			22041: outdata = 32'd43495;
			22042: outdata = 32'd43494;
			22043: outdata = 32'd43493;
			22044: outdata = 32'd43492;
			22045: outdata = 32'd43491;
			22046: outdata = 32'd43490;
			22047: outdata = 32'd43489;
			22048: outdata = 32'd43488;
			22049: outdata = 32'd43487;
			22050: outdata = 32'd43486;
			22051: outdata = 32'd43485;
			22052: outdata = 32'd43484;
			22053: outdata = 32'd43483;
			22054: outdata = 32'd43482;
			22055: outdata = 32'd43481;
			22056: outdata = 32'd43480;
			22057: outdata = 32'd43479;
			22058: outdata = 32'd43478;
			22059: outdata = 32'd43477;
			22060: outdata = 32'd43476;
			22061: outdata = 32'd43475;
			22062: outdata = 32'd43474;
			22063: outdata = 32'd43473;
			22064: outdata = 32'd43472;
			22065: outdata = 32'd43471;
			22066: outdata = 32'd43470;
			22067: outdata = 32'd43469;
			22068: outdata = 32'd43468;
			22069: outdata = 32'd43467;
			22070: outdata = 32'd43466;
			22071: outdata = 32'd43465;
			22072: outdata = 32'd43464;
			22073: outdata = 32'd43463;
			22074: outdata = 32'd43462;
			22075: outdata = 32'd43461;
			22076: outdata = 32'd43460;
			22077: outdata = 32'd43459;
			22078: outdata = 32'd43458;
			22079: outdata = 32'd43457;
			22080: outdata = 32'd43456;
			22081: outdata = 32'd43455;
			22082: outdata = 32'd43454;
			22083: outdata = 32'd43453;
			22084: outdata = 32'd43452;
			22085: outdata = 32'd43451;
			22086: outdata = 32'd43450;
			22087: outdata = 32'd43449;
			22088: outdata = 32'd43448;
			22089: outdata = 32'd43447;
			22090: outdata = 32'd43446;
			22091: outdata = 32'd43445;
			22092: outdata = 32'd43444;
			22093: outdata = 32'd43443;
			22094: outdata = 32'd43442;
			22095: outdata = 32'd43441;
			22096: outdata = 32'd43440;
			22097: outdata = 32'd43439;
			22098: outdata = 32'd43438;
			22099: outdata = 32'd43437;
			22100: outdata = 32'd43436;
			22101: outdata = 32'd43435;
			22102: outdata = 32'd43434;
			22103: outdata = 32'd43433;
			22104: outdata = 32'd43432;
			22105: outdata = 32'd43431;
			22106: outdata = 32'd43430;
			22107: outdata = 32'd43429;
			22108: outdata = 32'd43428;
			22109: outdata = 32'd43427;
			22110: outdata = 32'd43426;
			22111: outdata = 32'd43425;
			22112: outdata = 32'd43424;
			22113: outdata = 32'd43423;
			22114: outdata = 32'd43422;
			22115: outdata = 32'd43421;
			22116: outdata = 32'd43420;
			22117: outdata = 32'd43419;
			22118: outdata = 32'd43418;
			22119: outdata = 32'd43417;
			22120: outdata = 32'd43416;
			22121: outdata = 32'd43415;
			22122: outdata = 32'd43414;
			22123: outdata = 32'd43413;
			22124: outdata = 32'd43412;
			22125: outdata = 32'd43411;
			22126: outdata = 32'd43410;
			22127: outdata = 32'd43409;
			22128: outdata = 32'd43408;
			22129: outdata = 32'd43407;
			22130: outdata = 32'd43406;
			22131: outdata = 32'd43405;
			22132: outdata = 32'd43404;
			22133: outdata = 32'd43403;
			22134: outdata = 32'd43402;
			22135: outdata = 32'd43401;
			22136: outdata = 32'd43400;
			22137: outdata = 32'd43399;
			22138: outdata = 32'd43398;
			22139: outdata = 32'd43397;
			22140: outdata = 32'd43396;
			22141: outdata = 32'd43395;
			22142: outdata = 32'd43394;
			22143: outdata = 32'd43393;
			22144: outdata = 32'd43392;
			22145: outdata = 32'd43391;
			22146: outdata = 32'd43390;
			22147: outdata = 32'd43389;
			22148: outdata = 32'd43388;
			22149: outdata = 32'd43387;
			22150: outdata = 32'd43386;
			22151: outdata = 32'd43385;
			22152: outdata = 32'd43384;
			22153: outdata = 32'd43383;
			22154: outdata = 32'd43382;
			22155: outdata = 32'd43381;
			22156: outdata = 32'd43380;
			22157: outdata = 32'd43379;
			22158: outdata = 32'd43378;
			22159: outdata = 32'd43377;
			22160: outdata = 32'd43376;
			22161: outdata = 32'd43375;
			22162: outdata = 32'd43374;
			22163: outdata = 32'd43373;
			22164: outdata = 32'd43372;
			22165: outdata = 32'd43371;
			22166: outdata = 32'd43370;
			22167: outdata = 32'd43369;
			22168: outdata = 32'd43368;
			22169: outdata = 32'd43367;
			22170: outdata = 32'd43366;
			22171: outdata = 32'd43365;
			22172: outdata = 32'd43364;
			22173: outdata = 32'd43363;
			22174: outdata = 32'd43362;
			22175: outdata = 32'd43361;
			22176: outdata = 32'd43360;
			22177: outdata = 32'd43359;
			22178: outdata = 32'd43358;
			22179: outdata = 32'd43357;
			22180: outdata = 32'd43356;
			22181: outdata = 32'd43355;
			22182: outdata = 32'd43354;
			22183: outdata = 32'd43353;
			22184: outdata = 32'd43352;
			22185: outdata = 32'd43351;
			22186: outdata = 32'd43350;
			22187: outdata = 32'd43349;
			22188: outdata = 32'd43348;
			22189: outdata = 32'd43347;
			22190: outdata = 32'd43346;
			22191: outdata = 32'd43345;
			22192: outdata = 32'd43344;
			22193: outdata = 32'd43343;
			22194: outdata = 32'd43342;
			22195: outdata = 32'd43341;
			22196: outdata = 32'd43340;
			22197: outdata = 32'd43339;
			22198: outdata = 32'd43338;
			22199: outdata = 32'd43337;
			22200: outdata = 32'd43336;
			22201: outdata = 32'd43335;
			22202: outdata = 32'd43334;
			22203: outdata = 32'd43333;
			22204: outdata = 32'd43332;
			22205: outdata = 32'd43331;
			22206: outdata = 32'd43330;
			22207: outdata = 32'd43329;
			22208: outdata = 32'd43328;
			22209: outdata = 32'd43327;
			22210: outdata = 32'd43326;
			22211: outdata = 32'd43325;
			22212: outdata = 32'd43324;
			22213: outdata = 32'd43323;
			22214: outdata = 32'd43322;
			22215: outdata = 32'd43321;
			22216: outdata = 32'd43320;
			22217: outdata = 32'd43319;
			22218: outdata = 32'd43318;
			22219: outdata = 32'd43317;
			22220: outdata = 32'd43316;
			22221: outdata = 32'd43315;
			22222: outdata = 32'd43314;
			22223: outdata = 32'd43313;
			22224: outdata = 32'd43312;
			22225: outdata = 32'd43311;
			22226: outdata = 32'd43310;
			22227: outdata = 32'd43309;
			22228: outdata = 32'd43308;
			22229: outdata = 32'd43307;
			22230: outdata = 32'd43306;
			22231: outdata = 32'd43305;
			22232: outdata = 32'd43304;
			22233: outdata = 32'd43303;
			22234: outdata = 32'd43302;
			22235: outdata = 32'd43301;
			22236: outdata = 32'd43300;
			22237: outdata = 32'd43299;
			22238: outdata = 32'd43298;
			22239: outdata = 32'd43297;
			22240: outdata = 32'd43296;
			22241: outdata = 32'd43295;
			22242: outdata = 32'd43294;
			22243: outdata = 32'd43293;
			22244: outdata = 32'd43292;
			22245: outdata = 32'd43291;
			22246: outdata = 32'd43290;
			22247: outdata = 32'd43289;
			22248: outdata = 32'd43288;
			22249: outdata = 32'd43287;
			22250: outdata = 32'd43286;
			22251: outdata = 32'd43285;
			22252: outdata = 32'd43284;
			22253: outdata = 32'd43283;
			22254: outdata = 32'd43282;
			22255: outdata = 32'd43281;
			22256: outdata = 32'd43280;
			22257: outdata = 32'd43279;
			22258: outdata = 32'd43278;
			22259: outdata = 32'd43277;
			22260: outdata = 32'd43276;
			22261: outdata = 32'd43275;
			22262: outdata = 32'd43274;
			22263: outdata = 32'd43273;
			22264: outdata = 32'd43272;
			22265: outdata = 32'd43271;
			22266: outdata = 32'd43270;
			22267: outdata = 32'd43269;
			22268: outdata = 32'd43268;
			22269: outdata = 32'd43267;
			22270: outdata = 32'd43266;
			22271: outdata = 32'd43265;
			22272: outdata = 32'd43264;
			22273: outdata = 32'd43263;
			22274: outdata = 32'd43262;
			22275: outdata = 32'd43261;
			22276: outdata = 32'd43260;
			22277: outdata = 32'd43259;
			22278: outdata = 32'd43258;
			22279: outdata = 32'd43257;
			22280: outdata = 32'd43256;
			22281: outdata = 32'd43255;
			22282: outdata = 32'd43254;
			22283: outdata = 32'd43253;
			22284: outdata = 32'd43252;
			22285: outdata = 32'd43251;
			22286: outdata = 32'd43250;
			22287: outdata = 32'd43249;
			22288: outdata = 32'd43248;
			22289: outdata = 32'd43247;
			22290: outdata = 32'd43246;
			22291: outdata = 32'd43245;
			22292: outdata = 32'd43244;
			22293: outdata = 32'd43243;
			22294: outdata = 32'd43242;
			22295: outdata = 32'd43241;
			22296: outdata = 32'd43240;
			22297: outdata = 32'd43239;
			22298: outdata = 32'd43238;
			22299: outdata = 32'd43237;
			22300: outdata = 32'd43236;
			22301: outdata = 32'd43235;
			22302: outdata = 32'd43234;
			22303: outdata = 32'd43233;
			22304: outdata = 32'd43232;
			22305: outdata = 32'd43231;
			22306: outdata = 32'd43230;
			22307: outdata = 32'd43229;
			22308: outdata = 32'd43228;
			22309: outdata = 32'd43227;
			22310: outdata = 32'd43226;
			22311: outdata = 32'd43225;
			22312: outdata = 32'd43224;
			22313: outdata = 32'd43223;
			22314: outdata = 32'd43222;
			22315: outdata = 32'd43221;
			22316: outdata = 32'd43220;
			22317: outdata = 32'd43219;
			22318: outdata = 32'd43218;
			22319: outdata = 32'd43217;
			22320: outdata = 32'd43216;
			22321: outdata = 32'd43215;
			22322: outdata = 32'd43214;
			22323: outdata = 32'd43213;
			22324: outdata = 32'd43212;
			22325: outdata = 32'd43211;
			22326: outdata = 32'd43210;
			22327: outdata = 32'd43209;
			22328: outdata = 32'd43208;
			22329: outdata = 32'd43207;
			22330: outdata = 32'd43206;
			22331: outdata = 32'd43205;
			22332: outdata = 32'd43204;
			22333: outdata = 32'd43203;
			22334: outdata = 32'd43202;
			22335: outdata = 32'd43201;
			22336: outdata = 32'd43200;
			22337: outdata = 32'd43199;
			22338: outdata = 32'd43198;
			22339: outdata = 32'd43197;
			22340: outdata = 32'd43196;
			22341: outdata = 32'd43195;
			22342: outdata = 32'd43194;
			22343: outdata = 32'd43193;
			22344: outdata = 32'd43192;
			22345: outdata = 32'd43191;
			22346: outdata = 32'd43190;
			22347: outdata = 32'd43189;
			22348: outdata = 32'd43188;
			22349: outdata = 32'd43187;
			22350: outdata = 32'd43186;
			22351: outdata = 32'd43185;
			22352: outdata = 32'd43184;
			22353: outdata = 32'd43183;
			22354: outdata = 32'd43182;
			22355: outdata = 32'd43181;
			22356: outdata = 32'd43180;
			22357: outdata = 32'd43179;
			22358: outdata = 32'd43178;
			22359: outdata = 32'd43177;
			22360: outdata = 32'd43176;
			22361: outdata = 32'd43175;
			22362: outdata = 32'd43174;
			22363: outdata = 32'd43173;
			22364: outdata = 32'd43172;
			22365: outdata = 32'd43171;
			22366: outdata = 32'd43170;
			22367: outdata = 32'd43169;
			22368: outdata = 32'd43168;
			22369: outdata = 32'd43167;
			22370: outdata = 32'd43166;
			22371: outdata = 32'd43165;
			22372: outdata = 32'd43164;
			22373: outdata = 32'd43163;
			22374: outdata = 32'd43162;
			22375: outdata = 32'd43161;
			22376: outdata = 32'd43160;
			22377: outdata = 32'd43159;
			22378: outdata = 32'd43158;
			22379: outdata = 32'd43157;
			22380: outdata = 32'd43156;
			22381: outdata = 32'd43155;
			22382: outdata = 32'd43154;
			22383: outdata = 32'd43153;
			22384: outdata = 32'd43152;
			22385: outdata = 32'd43151;
			22386: outdata = 32'd43150;
			22387: outdata = 32'd43149;
			22388: outdata = 32'd43148;
			22389: outdata = 32'd43147;
			22390: outdata = 32'd43146;
			22391: outdata = 32'd43145;
			22392: outdata = 32'd43144;
			22393: outdata = 32'd43143;
			22394: outdata = 32'd43142;
			22395: outdata = 32'd43141;
			22396: outdata = 32'd43140;
			22397: outdata = 32'd43139;
			22398: outdata = 32'd43138;
			22399: outdata = 32'd43137;
			22400: outdata = 32'd43136;
			22401: outdata = 32'd43135;
			22402: outdata = 32'd43134;
			22403: outdata = 32'd43133;
			22404: outdata = 32'd43132;
			22405: outdata = 32'd43131;
			22406: outdata = 32'd43130;
			22407: outdata = 32'd43129;
			22408: outdata = 32'd43128;
			22409: outdata = 32'd43127;
			22410: outdata = 32'd43126;
			22411: outdata = 32'd43125;
			22412: outdata = 32'd43124;
			22413: outdata = 32'd43123;
			22414: outdata = 32'd43122;
			22415: outdata = 32'd43121;
			22416: outdata = 32'd43120;
			22417: outdata = 32'd43119;
			22418: outdata = 32'd43118;
			22419: outdata = 32'd43117;
			22420: outdata = 32'd43116;
			22421: outdata = 32'd43115;
			22422: outdata = 32'd43114;
			22423: outdata = 32'd43113;
			22424: outdata = 32'd43112;
			22425: outdata = 32'd43111;
			22426: outdata = 32'd43110;
			22427: outdata = 32'd43109;
			22428: outdata = 32'd43108;
			22429: outdata = 32'd43107;
			22430: outdata = 32'd43106;
			22431: outdata = 32'd43105;
			22432: outdata = 32'd43104;
			22433: outdata = 32'd43103;
			22434: outdata = 32'd43102;
			22435: outdata = 32'd43101;
			22436: outdata = 32'd43100;
			22437: outdata = 32'd43099;
			22438: outdata = 32'd43098;
			22439: outdata = 32'd43097;
			22440: outdata = 32'd43096;
			22441: outdata = 32'd43095;
			22442: outdata = 32'd43094;
			22443: outdata = 32'd43093;
			22444: outdata = 32'd43092;
			22445: outdata = 32'd43091;
			22446: outdata = 32'd43090;
			22447: outdata = 32'd43089;
			22448: outdata = 32'd43088;
			22449: outdata = 32'd43087;
			22450: outdata = 32'd43086;
			22451: outdata = 32'd43085;
			22452: outdata = 32'd43084;
			22453: outdata = 32'd43083;
			22454: outdata = 32'd43082;
			22455: outdata = 32'd43081;
			22456: outdata = 32'd43080;
			22457: outdata = 32'd43079;
			22458: outdata = 32'd43078;
			22459: outdata = 32'd43077;
			22460: outdata = 32'd43076;
			22461: outdata = 32'd43075;
			22462: outdata = 32'd43074;
			22463: outdata = 32'd43073;
			22464: outdata = 32'd43072;
			22465: outdata = 32'd43071;
			22466: outdata = 32'd43070;
			22467: outdata = 32'd43069;
			22468: outdata = 32'd43068;
			22469: outdata = 32'd43067;
			22470: outdata = 32'd43066;
			22471: outdata = 32'd43065;
			22472: outdata = 32'd43064;
			22473: outdata = 32'd43063;
			22474: outdata = 32'd43062;
			22475: outdata = 32'd43061;
			22476: outdata = 32'd43060;
			22477: outdata = 32'd43059;
			22478: outdata = 32'd43058;
			22479: outdata = 32'd43057;
			22480: outdata = 32'd43056;
			22481: outdata = 32'd43055;
			22482: outdata = 32'd43054;
			22483: outdata = 32'd43053;
			22484: outdata = 32'd43052;
			22485: outdata = 32'd43051;
			22486: outdata = 32'd43050;
			22487: outdata = 32'd43049;
			22488: outdata = 32'd43048;
			22489: outdata = 32'd43047;
			22490: outdata = 32'd43046;
			22491: outdata = 32'd43045;
			22492: outdata = 32'd43044;
			22493: outdata = 32'd43043;
			22494: outdata = 32'd43042;
			22495: outdata = 32'd43041;
			22496: outdata = 32'd43040;
			22497: outdata = 32'd43039;
			22498: outdata = 32'd43038;
			22499: outdata = 32'd43037;
			22500: outdata = 32'd43036;
			22501: outdata = 32'd43035;
			22502: outdata = 32'd43034;
			22503: outdata = 32'd43033;
			22504: outdata = 32'd43032;
			22505: outdata = 32'd43031;
			22506: outdata = 32'd43030;
			22507: outdata = 32'd43029;
			22508: outdata = 32'd43028;
			22509: outdata = 32'd43027;
			22510: outdata = 32'd43026;
			22511: outdata = 32'd43025;
			22512: outdata = 32'd43024;
			22513: outdata = 32'd43023;
			22514: outdata = 32'd43022;
			22515: outdata = 32'd43021;
			22516: outdata = 32'd43020;
			22517: outdata = 32'd43019;
			22518: outdata = 32'd43018;
			22519: outdata = 32'd43017;
			22520: outdata = 32'd43016;
			22521: outdata = 32'd43015;
			22522: outdata = 32'd43014;
			22523: outdata = 32'd43013;
			22524: outdata = 32'd43012;
			22525: outdata = 32'd43011;
			22526: outdata = 32'd43010;
			22527: outdata = 32'd43009;
			22528: outdata = 32'd43008;
			22529: outdata = 32'd43007;
			22530: outdata = 32'd43006;
			22531: outdata = 32'd43005;
			22532: outdata = 32'd43004;
			22533: outdata = 32'd43003;
			22534: outdata = 32'd43002;
			22535: outdata = 32'd43001;
			22536: outdata = 32'd43000;
			22537: outdata = 32'd42999;
			22538: outdata = 32'd42998;
			22539: outdata = 32'd42997;
			22540: outdata = 32'd42996;
			22541: outdata = 32'd42995;
			22542: outdata = 32'd42994;
			22543: outdata = 32'd42993;
			22544: outdata = 32'd42992;
			22545: outdata = 32'd42991;
			22546: outdata = 32'd42990;
			22547: outdata = 32'd42989;
			22548: outdata = 32'd42988;
			22549: outdata = 32'd42987;
			22550: outdata = 32'd42986;
			22551: outdata = 32'd42985;
			22552: outdata = 32'd42984;
			22553: outdata = 32'd42983;
			22554: outdata = 32'd42982;
			22555: outdata = 32'd42981;
			22556: outdata = 32'd42980;
			22557: outdata = 32'd42979;
			22558: outdata = 32'd42978;
			22559: outdata = 32'd42977;
			22560: outdata = 32'd42976;
			22561: outdata = 32'd42975;
			22562: outdata = 32'd42974;
			22563: outdata = 32'd42973;
			22564: outdata = 32'd42972;
			22565: outdata = 32'd42971;
			22566: outdata = 32'd42970;
			22567: outdata = 32'd42969;
			22568: outdata = 32'd42968;
			22569: outdata = 32'd42967;
			22570: outdata = 32'd42966;
			22571: outdata = 32'd42965;
			22572: outdata = 32'd42964;
			22573: outdata = 32'd42963;
			22574: outdata = 32'd42962;
			22575: outdata = 32'd42961;
			22576: outdata = 32'd42960;
			22577: outdata = 32'd42959;
			22578: outdata = 32'd42958;
			22579: outdata = 32'd42957;
			22580: outdata = 32'd42956;
			22581: outdata = 32'd42955;
			22582: outdata = 32'd42954;
			22583: outdata = 32'd42953;
			22584: outdata = 32'd42952;
			22585: outdata = 32'd42951;
			22586: outdata = 32'd42950;
			22587: outdata = 32'd42949;
			22588: outdata = 32'd42948;
			22589: outdata = 32'd42947;
			22590: outdata = 32'd42946;
			22591: outdata = 32'd42945;
			22592: outdata = 32'd42944;
			22593: outdata = 32'd42943;
			22594: outdata = 32'd42942;
			22595: outdata = 32'd42941;
			22596: outdata = 32'd42940;
			22597: outdata = 32'd42939;
			22598: outdata = 32'd42938;
			22599: outdata = 32'd42937;
			22600: outdata = 32'd42936;
			22601: outdata = 32'd42935;
			22602: outdata = 32'd42934;
			22603: outdata = 32'd42933;
			22604: outdata = 32'd42932;
			22605: outdata = 32'd42931;
			22606: outdata = 32'd42930;
			22607: outdata = 32'd42929;
			22608: outdata = 32'd42928;
			22609: outdata = 32'd42927;
			22610: outdata = 32'd42926;
			22611: outdata = 32'd42925;
			22612: outdata = 32'd42924;
			22613: outdata = 32'd42923;
			22614: outdata = 32'd42922;
			22615: outdata = 32'd42921;
			22616: outdata = 32'd42920;
			22617: outdata = 32'd42919;
			22618: outdata = 32'd42918;
			22619: outdata = 32'd42917;
			22620: outdata = 32'd42916;
			22621: outdata = 32'd42915;
			22622: outdata = 32'd42914;
			22623: outdata = 32'd42913;
			22624: outdata = 32'd42912;
			22625: outdata = 32'd42911;
			22626: outdata = 32'd42910;
			22627: outdata = 32'd42909;
			22628: outdata = 32'd42908;
			22629: outdata = 32'd42907;
			22630: outdata = 32'd42906;
			22631: outdata = 32'd42905;
			22632: outdata = 32'd42904;
			22633: outdata = 32'd42903;
			22634: outdata = 32'd42902;
			22635: outdata = 32'd42901;
			22636: outdata = 32'd42900;
			22637: outdata = 32'd42899;
			22638: outdata = 32'd42898;
			22639: outdata = 32'd42897;
			22640: outdata = 32'd42896;
			22641: outdata = 32'd42895;
			22642: outdata = 32'd42894;
			22643: outdata = 32'd42893;
			22644: outdata = 32'd42892;
			22645: outdata = 32'd42891;
			22646: outdata = 32'd42890;
			22647: outdata = 32'd42889;
			22648: outdata = 32'd42888;
			22649: outdata = 32'd42887;
			22650: outdata = 32'd42886;
			22651: outdata = 32'd42885;
			22652: outdata = 32'd42884;
			22653: outdata = 32'd42883;
			22654: outdata = 32'd42882;
			22655: outdata = 32'd42881;
			22656: outdata = 32'd42880;
			22657: outdata = 32'd42879;
			22658: outdata = 32'd42878;
			22659: outdata = 32'd42877;
			22660: outdata = 32'd42876;
			22661: outdata = 32'd42875;
			22662: outdata = 32'd42874;
			22663: outdata = 32'd42873;
			22664: outdata = 32'd42872;
			22665: outdata = 32'd42871;
			22666: outdata = 32'd42870;
			22667: outdata = 32'd42869;
			22668: outdata = 32'd42868;
			22669: outdata = 32'd42867;
			22670: outdata = 32'd42866;
			22671: outdata = 32'd42865;
			22672: outdata = 32'd42864;
			22673: outdata = 32'd42863;
			22674: outdata = 32'd42862;
			22675: outdata = 32'd42861;
			22676: outdata = 32'd42860;
			22677: outdata = 32'd42859;
			22678: outdata = 32'd42858;
			22679: outdata = 32'd42857;
			22680: outdata = 32'd42856;
			22681: outdata = 32'd42855;
			22682: outdata = 32'd42854;
			22683: outdata = 32'd42853;
			22684: outdata = 32'd42852;
			22685: outdata = 32'd42851;
			22686: outdata = 32'd42850;
			22687: outdata = 32'd42849;
			22688: outdata = 32'd42848;
			22689: outdata = 32'd42847;
			22690: outdata = 32'd42846;
			22691: outdata = 32'd42845;
			22692: outdata = 32'd42844;
			22693: outdata = 32'd42843;
			22694: outdata = 32'd42842;
			22695: outdata = 32'd42841;
			22696: outdata = 32'd42840;
			22697: outdata = 32'd42839;
			22698: outdata = 32'd42838;
			22699: outdata = 32'd42837;
			22700: outdata = 32'd42836;
			22701: outdata = 32'd42835;
			22702: outdata = 32'd42834;
			22703: outdata = 32'd42833;
			22704: outdata = 32'd42832;
			22705: outdata = 32'd42831;
			22706: outdata = 32'd42830;
			22707: outdata = 32'd42829;
			22708: outdata = 32'd42828;
			22709: outdata = 32'd42827;
			22710: outdata = 32'd42826;
			22711: outdata = 32'd42825;
			22712: outdata = 32'd42824;
			22713: outdata = 32'd42823;
			22714: outdata = 32'd42822;
			22715: outdata = 32'd42821;
			22716: outdata = 32'd42820;
			22717: outdata = 32'd42819;
			22718: outdata = 32'd42818;
			22719: outdata = 32'd42817;
			22720: outdata = 32'd42816;
			22721: outdata = 32'd42815;
			22722: outdata = 32'd42814;
			22723: outdata = 32'd42813;
			22724: outdata = 32'd42812;
			22725: outdata = 32'd42811;
			22726: outdata = 32'd42810;
			22727: outdata = 32'd42809;
			22728: outdata = 32'd42808;
			22729: outdata = 32'd42807;
			22730: outdata = 32'd42806;
			22731: outdata = 32'd42805;
			22732: outdata = 32'd42804;
			22733: outdata = 32'd42803;
			22734: outdata = 32'd42802;
			22735: outdata = 32'd42801;
			22736: outdata = 32'd42800;
			22737: outdata = 32'd42799;
			22738: outdata = 32'd42798;
			22739: outdata = 32'd42797;
			22740: outdata = 32'd42796;
			22741: outdata = 32'd42795;
			22742: outdata = 32'd42794;
			22743: outdata = 32'd42793;
			22744: outdata = 32'd42792;
			22745: outdata = 32'd42791;
			22746: outdata = 32'd42790;
			22747: outdata = 32'd42789;
			22748: outdata = 32'd42788;
			22749: outdata = 32'd42787;
			22750: outdata = 32'd42786;
			22751: outdata = 32'd42785;
			22752: outdata = 32'd42784;
			22753: outdata = 32'd42783;
			22754: outdata = 32'd42782;
			22755: outdata = 32'd42781;
			22756: outdata = 32'd42780;
			22757: outdata = 32'd42779;
			22758: outdata = 32'd42778;
			22759: outdata = 32'd42777;
			22760: outdata = 32'd42776;
			22761: outdata = 32'd42775;
			22762: outdata = 32'd42774;
			22763: outdata = 32'd42773;
			22764: outdata = 32'd42772;
			22765: outdata = 32'd42771;
			22766: outdata = 32'd42770;
			22767: outdata = 32'd42769;
			22768: outdata = 32'd42768;
			22769: outdata = 32'd42767;
			22770: outdata = 32'd42766;
			22771: outdata = 32'd42765;
			22772: outdata = 32'd42764;
			22773: outdata = 32'd42763;
			22774: outdata = 32'd42762;
			22775: outdata = 32'd42761;
			22776: outdata = 32'd42760;
			22777: outdata = 32'd42759;
			22778: outdata = 32'd42758;
			22779: outdata = 32'd42757;
			22780: outdata = 32'd42756;
			22781: outdata = 32'd42755;
			22782: outdata = 32'd42754;
			22783: outdata = 32'd42753;
			22784: outdata = 32'd42752;
			22785: outdata = 32'd42751;
			22786: outdata = 32'd42750;
			22787: outdata = 32'd42749;
			22788: outdata = 32'd42748;
			22789: outdata = 32'd42747;
			22790: outdata = 32'd42746;
			22791: outdata = 32'd42745;
			22792: outdata = 32'd42744;
			22793: outdata = 32'd42743;
			22794: outdata = 32'd42742;
			22795: outdata = 32'd42741;
			22796: outdata = 32'd42740;
			22797: outdata = 32'd42739;
			22798: outdata = 32'd42738;
			22799: outdata = 32'd42737;
			22800: outdata = 32'd42736;
			22801: outdata = 32'd42735;
			22802: outdata = 32'd42734;
			22803: outdata = 32'd42733;
			22804: outdata = 32'd42732;
			22805: outdata = 32'd42731;
			22806: outdata = 32'd42730;
			22807: outdata = 32'd42729;
			22808: outdata = 32'd42728;
			22809: outdata = 32'd42727;
			22810: outdata = 32'd42726;
			22811: outdata = 32'd42725;
			22812: outdata = 32'd42724;
			22813: outdata = 32'd42723;
			22814: outdata = 32'd42722;
			22815: outdata = 32'd42721;
			22816: outdata = 32'd42720;
			22817: outdata = 32'd42719;
			22818: outdata = 32'd42718;
			22819: outdata = 32'd42717;
			22820: outdata = 32'd42716;
			22821: outdata = 32'd42715;
			22822: outdata = 32'd42714;
			22823: outdata = 32'd42713;
			22824: outdata = 32'd42712;
			22825: outdata = 32'd42711;
			22826: outdata = 32'd42710;
			22827: outdata = 32'd42709;
			22828: outdata = 32'd42708;
			22829: outdata = 32'd42707;
			22830: outdata = 32'd42706;
			22831: outdata = 32'd42705;
			22832: outdata = 32'd42704;
			22833: outdata = 32'd42703;
			22834: outdata = 32'd42702;
			22835: outdata = 32'd42701;
			22836: outdata = 32'd42700;
			22837: outdata = 32'd42699;
			22838: outdata = 32'd42698;
			22839: outdata = 32'd42697;
			22840: outdata = 32'd42696;
			22841: outdata = 32'd42695;
			22842: outdata = 32'd42694;
			22843: outdata = 32'd42693;
			22844: outdata = 32'd42692;
			22845: outdata = 32'd42691;
			22846: outdata = 32'd42690;
			22847: outdata = 32'd42689;
			22848: outdata = 32'd42688;
			22849: outdata = 32'd42687;
			22850: outdata = 32'd42686;
			22851: outdata = 32'd42685;
			22852: outdata = 32'd42684;
			22853: outdata = 32'd42683;
			22854: outdata = 32'd42682;
			22855: outdata = 32'd42681;
			22856: outdata = 32'd42680;
			22857: outdata = 32'd42679;
			22858: outdata = 32'd42678;
			22859: outdata = 32'd42677;
			22860: outdata = 32'd42676;
			22861: outdata = 32'd42675;
			22862: outdata = 32'd42674;
			22863: outdata = 32'd42673;
			22864: outdata = 32'd42672;
			22865: outdata = 32'd42671;
			22866: outdata = 32'd42670;
			22867: outdata = 32'd42669;
			22868: outdata = 32'd42668;
			22869: outdata = 32'd42667;
			22870: outdata = 32'd42666;
			22871: outdata = 32'd42665;
			22872: outdata = 32'd42664;
			22873: outdata = 32'd42663;
			22874: outdata = 32'd42662;
			22875: outdata = 32'd42661;
			22876: outdata = 32'd42660;
			22877: outdata = 32'd42659;
			22878: outdata = 32'd42658;
			22879: outdata = 32'd42657;
			22880: outdata = 32'd42656;
			22881: outdata = 32'd42655;
			22882: outdata = 32'd42654;
			22883: outdata = 32'd42653;
			22884: outdata = 32'd42652;
			22885: outdata = 32'd42651;
			22886: outdata = 32'd42650;
			22887: outdata = 32'd42649;
			22888: outdata = 32'd42648;
			22889: outdata = 32'd42647;
			22890: outdata = 32'd42646;
			22891: outdata = 32'd42645;
			22892: outdata = 32'd42644;
			22893: outdata = 32'd42643;
			22894: outdata = 32'd42642;
			22895: outdata = 32'd42641;
			22896: outdata = 32'd42640;
			22897: outdata = 32'd42639;
			22898: outdata = 32'd42638;
			22899: outdata = 32'd42637;
			22900: outdata = 32'd42636;
			22901: outdata = 32'd42635;
			22902: outdata = 32'd42634;
			22903: outdata = 32'd42633;
			22904: outdata = 32'd42632;
			22905: outdata = 32'd42631;
			22906: outdata = 32'd42630;
			22907: outdata = 32'd42629;
			22908: outdata = 32'd42628;
			22909: outdata = 32'd42627;
			22910: outdata = 32'd42626;
			22911: outdata = 32'd42625;
			22912: outdata = 32'd42624;
			22913: outdata = 32'd42623;
			22914: outdata = 32'd42622;
			22915: outdata = 32'd42621;
			22916: outdata = 32'd42620;
			22917: outdata = 32'd42619;
			22918: outdata = 32'd42618;
			22919: outdata = 32'd42617;
			22920: outdata = 32'd42616;
			22921: outdata = 32'd42615;
			22922: outdata = 32'd42614;
			22923: outdata = 32'd42613;
			22924: outdata = 32'd42612;
			22925: outdata = 32'd42611;
			22926: outdata = 32'd42610;
			22927: outdata = 32'd42609;
			22928: outdata = 32'd42608;
			22929: outdata = 32'd42607;
			22930: outdata = 32'd42606;
			22931: outdata = 32'd42605;
			22932: outdata = 32'd42604;
			22933: outdata = 32'd42603;
			22934: outdata = 32'd42602;
			22935: outdata = 32'd42601;
			22936: outdata = 32'd42600;
			22937: outdata = 32'd42599;
			22938: outdata = 32'd42598;
			22939: outdata = 32'd42597;
			22940: outdata = 32'd42596;
			22941: outdata = 32'd42595;
			22942: outdata = 32'd42594;
			22943: outdata = 32'd42593;
			22944: outdata = 32'd42592;
			22945: outdata = 32'd42591;
			22946: outdata = 32'd42590;
			22947: outdata = 32'd42589;
			22948: outdata = 32'd42588;
			22949: outdata = 32'd42587;
			22950: outdata = 32'd42586;
			22951: outdata = 32'd42585;
			22952: outdata = 32'd42584;
			22953: outdata = 32'd42583;
			22954: outdata = 32'd42582;
			22955: outdata = 32'd42581;
			22956: outdata = 32'd42580;
			22957: outdata = 32'd42579;
			22958: outdata = 32'd42578;
			22959: outdata = 32'd42577;
			22960: outdata = 32'd42576;
			22961: outdata = 32'd42575;
			22962: outdata = 32'd42574;
			22963: outdata = 32'd42573;
			22964: outdata = 32'd42572;
			22965: outdata = 32'd42571;
			22966: outdata = 32'd42570;
			22967: outdata = 32'd42569;
			22968: outdata = 32'd42568;
			22969: outdata = 32'd42567;
			22970: outdata = 32'd42566;
			22971: outdata = 32'd42565;
			22972: outdata = 32'd42564;
			22973: outdata = 32'd42563;
			22974: outdata = 32'd42562;
			22975: outdata = 32'd42561;
			22976: outdata = 32'd42560;
			22977: outdata = 32'd42559;
			22978: outdata = 32'd42558;
			22979: outdata = 32'd42557;
			22980: outdata = 32'd42556;
			22981: outdata = 32'd42555;
			22982: outdata = 32'd42554;
			22983: outdata = 32'd42553;
			22984: outdata = 32'd42552;
			22985: outdata = 32'd42551;
			22986: outdata = 32'd42550;
			22987: outdata = 32'd42549;
			22988: outdata = 32'd42548;
			22989: outdata = 32'd42547;
			22990: outdata = 32'd42546;
			22991: outdata = 32'd42545;
			22992: outdata = 32'd42544;
			22993: outdata = 32'd42543;
			22994: outdata = 32'd42542;
			22995: outdata = 32'd42541;
			22996: outdata = 32'd42540;
			22997: outdata = 32'd42539;
			22998: outdata = 32'd42538;
			22999: outdata = 32'd42537;
			23000: outdata = 32'd42536;
			23001: outdata = 32'd42535;
			23002: outdata = 32'd42534;
			23003: outdata = 32'd42533;
			23004: outdata = 32'd42532;
			23005: outdata = 32'd42531;
			23006: outdata = 32'd42530;
			23007: outdata = 32'd42529;
			23008: outdata = 32'd42528;
			23009: outdata = 32'd42527;
			23010: outdata = 32'd42526;
			23011: outdata = 32'd42525;
			23012: outdata = 32'd42524;
			23013: outdata = 32'd42523;
			23014: outdata = 32'd42522;
			23015: outdata = 32'd42521;
			23016: outdata = 32'd42520;
			23017: outdata = 32'd42519;
			23018: outdata = 32'd42518;
			23019: outdata = 32'd42517;
			23020: outdata = 32'd42516;
			23021: outdata = 32'd42515;
			23022: outdata = 32'd42514;
			23023: outdata = 32'd42513;
			23024: outdata = 32'd42512;
			23025: outdata = 32'd42511;
			23026: outdata = 32'd42510;
			23027: outdata = 32'd42509;
			23028: outdata = 32'd42508;
			23029: outdata = 32'd42507;
			23030: outdata = 32'd42506;
			23031: outdata = 32'd42505;
			23032: outdata = 32'd42504;
			23033: outdata = 32'd42503;
			23034: outdata = 32'd42502;
			23035: outdata = 32'd42501;
			23036: outdata = 32'd42500;
			23037: outdata = 32'd42499;
			23038: outdata = 32'd42498;
			23039: outdata = 32'd42497;
			23040: outdata = 32'd42496;
			23041: outdata = 32'd42495;
			23042: outdata = 32'd42494;
			23043: outdata = 32'd42493;
			23044: outdata = 32'd42492;
			23045: outdata = 32'd42491;
			23046: outdata = 32'd42490;
			23047: outdata = 32'd42489;
			23048: outdata = 32'd42488;
			23049: outdata = 32'd42487;
			23050: outdata = 32'd42486;
			23051: outdata = 32'd42485;
			23052: outdata = 32'd42484;
			23053: outdata = 32'd42483;
			23054: outdata = 32'd42482;
			23055: outdata = 32'd42481;
			23056: outdata = 32'd42480;
			23057: outdata = 32'd42479;
			23058: outdata = 32'd42478;
			23059: outdata = 32'd42477;
			23060: outdata = 32'd42476;
			23061: outdata = 32'd42475;
			23062: outdata = 32'd42474;
			23063: outdata = 32'd42473;
			23064: outdata = 32'd42472;
			23065: outdata = 32'd42471;
			23066: outdata = 32'd42470;
			23067: outdata = 32'd42469;
			23068: outdata = 32'd42468;
			23069: outdata = 32'd42467;
			23070: outdata = 32'd42466;
			23071: outdata = 32'd42465;
			23072: outdata = 32'd42464;
			23073: outdata = 32'd42463;
			23074: outdata = 32'd42462;
			23075: outdata = 32'd42461;
			23076: outdata = 32'd42460;
			23077: outdata = 32'd42459;
			23078: outdata = 32'd42458;
			23079: outdata = 32'd42457;
			23080: outdata = 32'd42456;
			23081: outdata = 32'd42455;
			23082: outdata = 32'd42454;
			23083: outdata = 32'd42453;
			23084: outdata = 32'd42452;
			23085: outdata = 32'd42451;
			23086: outdata = 32'd42450;
			23087: outdata = 32'd42449;
			23088: outdata = 32'd42448;
			23089: outdata = 32'd42447;
			23090: outdata = 32'd42446;
			23091: outdata = 32'd42445;
			23092: outdata = 32'd42444;
			23093: outdata = 32'd42443;
			23094: outdata = 32'd42442;
			23095: outdata = 32'd42441;
			23096: outdata = 32'd42440;
			23097: outdata = 32'd42439;
			23098: outdata = 32'd42438;
			23099: outdata = 32'd42437;
			23100: outdata = 32'd42436;
			23101: outdata = 32'd42435;
			23102: outdata = 32'd42434;
			23103: outdata = 32'd42433;
			23104: outdata = 32'd42432;
			23105: outdata = 32'd42431;
			23106: outdata = 32'd42430;
			23107: outdata = 32'd42429;
			23108: outdata = 32'd42428;
			23109: outdata = 32'd42427;
			23110: outdata = 32'd42426;
			23111: outdata = 32'd42425;
			23112: outdata = 32'd42424;
			23113: outdata = 32'd42423;
			23114: outdata = 32'd42422;
			23115: outdata = 32'd42421;
			23116: outdata = 32'd42420;
			23117: outdata = 32'd42419;
			23118: outdata = 32'd42418;
			23119: outdata = 32'd42417;
			23120: outdata = 32'd42416;
			23121: outdata = 32'd42415;
			23122: outdata = 32'd42414;
			23123: outdata = 32'd42413;
			23124: outdata = 32'd42412;
			23125: outdata = 32'd42411;
			23126: outdata = 32'd42410;
			23127: outdata = 32'd42409;
			23128: outdata = 32'd42408;
			23129: outdata = 32'd42407;
			23130: outdata = 32'd42406;
			23131: outdata = 32'd42405;
			23132: outdata = 32'd42404;
			23133: outdata = 32'd42403;
			23134: outdata = 32'd42402;
			23135: outdata = 32'd42401;
			23136: outdata = 32'd42400;
			23137: outdata = 32'd42399;
			23138: outdata = 32'd42398;
			23139: outdata = 32'd42397;
			23140: outdata = 32'd42396;
			23141: outdata = 32'd42395;
			23142: outdata = 32'd42394;
			23143: outdata = 32'd42393;
			23144: outdata = 32'd42392;
			23145: outdata = 32'd42391;
			23146: outdata = 32'd42390;
			23147: outdata = 32'd42389;
			23148: outdata = 32'd42388;
			23149: outdata = 32'd42387;
			23150: outdata = 32'd42386;
			23151: outdata = 32'd42385;
			23152: outdata = 32'd42384;
			23153: outdata = 32'd42383;
			23154: outdata = 32'd42382;
			23155: outdata = 32'd42381;
			23156: outdata = 32'd42380;
			23157: outdata = 32'd42379;
			23158: outdata = 32'd42378;
			23159: outdata = 32'd42377;
			23160: outdata = 32'd42376;
			23161: outdata = 32'd42375;
			23162: outdata = 32'd42374;
			23163: outdata = 32'd42373;
			23164: outdata = 32'd42372;
			23165: outdata = 32'd42371;
			23166: outdata = 32'd42370;
			23167: outdata = 32'd42369;
			23168: outdata = 32'd42368;
			23169: outdata = 32'd42367;
			23170: outdata = 32'd42366;
			23171: outdata = 32'd42365;
			23172: outdata = 32'd42364;
			23173: outdata = 32'd42363;
			23174: outdata = 32'd42362;
			23175: outdata = 32'd42361;
			23176: outdata = 32'd42360;
			23177: outdata = 32'd42359;
			23178: outdata = 32'd42358;
			23179: outdata = 32'd42357;
			23180: outdata = 32'd42356;
			23181: outdata = 32'd42355;
			23182: outdata = 32'd42354;
			23183: outdata = 32'd42353;
			23184: outdata = 32'd42352;
			23185: outdata = 32'd42351;
			23186: outdata = 32'd42350;
			23187: outdata = 32'd42349;
			23188: outdata = 32'd42348;
			23189: outdata = 32'd42347;
			23190: outdata = 32'd42346;
			23191: outdata = 32'd42345;
			23192: outdata = 32'd42344;
			23193: outdata = 32'd42343;
			23194: outdata = 32'd42342;
			23195: outdata = 32'd42341;
			23196: outdata = 32'd42340;
			23197: outdata = 32'd42339;
			23198: outdata = 32'd42338;
			23199: outdata = 32'd42337;
			23200: outdata = 32'd42336;
			23201: outdata = 32'd42335;
			23202: outdata = 32'd42334;
			23203: outdata = 32'd42333;
			23204: outdata = 32'd42332;
			23205: outdata = 32'd42331;
			23206: outdata = 32'd42330;
			23207: outdata = 32'd42329;
			23208: outdata = 32'd42328;
			23209: outdata = 32'd42327;
			23210: outdata = 32'd42326;
			23211: outdata = 32'd42325;
			23212: outdata = 32'd42324;
			23213: outdata = 32'd42323;
			23214: outdata = 32'd42322;
			23215: outdata = 32'd42321;
			23216: outdata = 32'd42320;
			23217: outdata = 32'd42319;
			23218: outdata = 32'd42318;
			23219: outdata = 32'd42317;
			23220: outdata = 32'd42316;
			23221: outdata = 32'd42315;
			23222: outdata = 32'd42314;
			23223: outdata = 32'd42313;
			23224: outdata = 32'd42312;
			23225: outdata = 32'd42311;
			23226: outdata = 32'd42310;
			23227: outdata = 32'd42309;
			23228: outdata = 32'd42308;
			23229: outdata = 32'd42307;
			23230: outdata = 32'd42306;
			23231: outdata = 32'd42305;
			23232: outdata = 32'd42304;
			23233: outdata = 32'd42303;
			23234: outdata = 32'd42302;
			23235: outdata = 32'd42301;
			23236: outdata = 32'd42300;
			23237: outdata = 32'd42299;
			23238: outdata = 32'd42298;
			23239: outdata = 32'd42297;
			23240: outdata = 32'd42296;
			23241: outdata = 32'd42295;
			23242: outdata = 32'd42294;
			23243: outdata = 32'd42293;
			23244: outdata = 32'd42292;
			23245: outdata = 32'd42291;
			23246: outdata = 32'd42290;
			23247: outdata = 32'd42289;
			23248: outdata = 32'd42288;
			23249: outdata = 32'd42287;
			23250: outdata = 32'd42286;
			23251: outdata = 32'd42285;
			23252: outdata = 32'd42284;
			23253: outdata = 32'd42283;
			23254: outdata = 32'd42282;
			23255: outdata = 32'd42281;
			23256: outdata = 32'd42280;
			23257: outdata = 32'd42279;
			23258: outdata = 32'd42278;
			23259: outdata = 32'd42277;
			23260: outdata = 32'd42276;
			23261: outdata = 32'd42275;
			23262: outdata = 32'd42274;
			23263: outdata = 32'd42273;
			23264: outdata = 32'd42272;
			23265: outdata = 32'd42271;
			23266: outdata = 32'd42270;
			23267: outdata = 32'd42269;
			23268: outdata = 32'd42268;
			23269: outdata = 32'd42267;
			23270: outdata = 32'd42266;
			23271: outdata = 32'd42265;
			23272: outdata = 32'd42264;
			23273: outdata = 32'd42263;
			23274: outdata = 32'd42262;
			23275: outdata = 32'd42261;
			23276: outdata = 32'd42260;
			23277: outdata = 32'd42259;
			23278: outdata = 32'd42258;
			23279: outdata = 32'd42257;
			23280: outdata = 32'd42256;
			23281: outdata = 32'd42255;
			23282: outdata = 32'd42254;
			23283: outdata = 32'd42253;
			23284: outdata = 32'd42252;
			23285: outdata = 32'd42251;
			23286: outdata = 32'd42250;
			23287: outdata = 32'd42249;
			23288: outdata = 32'd42248;
			23289: outdata = 32'd42247;
			23290: outdata = 32'd42246;
			23291: outdata = 32'd42245;
			23292: outdata = 32'd42244;
			23293: outdata = 32'd42243;
			23294: outdata = 32'd42242;
			23295: outdata = 32'd42241;
			23296: outdata = 32'd42240;
			23297: outdata = 32'd42239;
			23298: outdata = 32'd42238;
			23299: outdata = 32'd42237;
			23300: outdata = 32'd42236;
			23301: outdata = 32'd42235;
			23302: outdata = 32'd42234;
			23303: outdata = 32'd42233;
			23304: outdata = 32'd42232;
			23305: outdata = 32'd42231;
			23306: outdata = 32'd42230;
			23307: outdata = 32'd42229;
			23308: outdata = 32'd42228;
			23309: outdata = 32'd42227;
			23310: outdata = 32'd42226;
			23311: outdata = 32'd42225;
			23312: outdata = 32'd42224;
			23313: outdata = 32'd42223;
			23314: outdata = 32'd42222;
			23315: outdata = 32'd42221;
			23316: outdata = 32'd42220;
			23317: outdata = 32'd42219;
			23318: outdata = 32'd42218;
			23319: outdata = 32'd42217;
			23320: outdata = 32'd42216;
			23321: outdata = 32'd42215;
			23322: outdata = 32'd42214;
			23323: outdata = 32'd42213;
			23324: outdata = 32'd42212;
			23325: outdata = 32'd42211;
			23326: outdata = 32'd42210;
			23327: outdata = 32'd42209;
			23328: outdata = 32'd42208;
			23329: outdata = 32'd42207;
			23330: outdata = 32'd42206;
			23331: outdata = 32'd42205;
			23332: outdata = 32'd42204;
			23333: outdata = 32'd42203;
			23334: outdata = 32'd42202;
			23335: outdata = 32'd42201;
			23336: outdata = 32'd42200;
			23337: outdata = 32'd42199;
			23338: outdata = 32'd42198;
			23339: outdata = 32'd42197;
			23340: outdata = 32'd42196;
			23341: outdata = 32'd42195;
			23342: outdata = 32'd42194;
			23343: outdata = 32'd42193;
			23344: outdata = 32'd42192;
			23345: outdata = 32'd42191;
			23346: outdata = 32'd42190;
			23347: outdata = 32'd42189;
			23348: outdata = 32'd42188;
			23349: outdata = 32'd42187;
			23350: outdata = 32'd42186;
			23351: outdata = 32'd42185;
			23352: outdata = 32'd42184;
			23353: outdata = 32'd42183;
			23354: outdata = 32'd42182;
			23355: outdata = 32'd42181;
			23356: outdata = 32'd42180;
			23357: outdata = 32'd42179;
			23358: outdata = 32'd42178;
			23359: outdata = 32'd42177;
			23360: outdata = 32'd42176;
			23361: outdata = 32'd42175;
			23362: outdata = 32'd42174;
			23363: outdata = 32'd42173;
			23364: outdata = 32'd42172;
			23365: outdata = 32'd42171;
			23366: outdata = 32'd42170;
			23367: outdata = 32'd42169;
			23368: outdata = 32'd42168;
			23369: outdata = 32'd42167;
			23370: outdata = 32'd42166;
			23371: outdata = 32'd42165;
			23372: outdata = 32'd42164;
			23373: outdata = 32'd42163;
			23374: outdata = 32'd42162;
			23375: outdata = 32'd42161;
			23376: outdata = 32'd42160;
			23377: outdata = 32'd42159;
			23378: outdata = 32'd42158;
			23379: outdata = 32'd42157;
			23380: outdata = 32'd42156;
			23381: outdata = 32'd42155;
			23382: outdata = 32'd42154;
			23383: outdata = 32'd42153;
			23384: outdata = 32'd42152;
			23385: outdata = 32'd42151;
			23386: outdata = 32'd42150;
			23387: outdata = 32'd42149;
			23388: outdata = 32'd42148;
			23389: outdata = 32'd42147;
			23390: outdata = 32'd42146;
			23391: outdata = 32'd42145;
			23392: outdata = 32'd42144;
			23393: outdata = 32'd42143;
			23394: outdata = 32'd42142;
			23395: outdata = 32'd42141;
			23396: outdata = 32'd42140;
			23397: outdata = 32'd42139;
			23398: outdata = 32'd42138;
			23399: outdata = 32'd42137;
			23400: outdata = 32'd42136;
			23401: outdata = 32'd42135;
			23402: outdata = 32'd42134;
			23403: outdata = 32'd42133;
			23404: outdata = 32'd42132;
			23405: outdata = 32'd42131;
			23406: outdata = 32'd42130;
			23407: outdata = 32'd42129;
			23408: outdata = 32'd42128;
			23409: outdata = 32'd42127;
			23410: outdata = 32'd42126;
			23411: outdata = 32'd42125;
			23412: outdata = 32'd42124;
			23413: outdata = 32'd42123;
			23414: outdata = 32'd42122;
			23415: outdata = 32'd42121;
			23416: outdata = 32'd42120;
			23417: outdata = 32'd42119;
			23418: outdata = 32'd42118;
			23419: outdata = 32'd42117;
			23420: outdata = 32'd42116;
			23421: outdata = 32'd42115;
			23422: outdata = 32'd42114;
			23423: outdata = 32'd42113;
			23424: outdata = 32'd42112;
			23425: outdata = 32'd42111;
			23426: outdata = 32'd42110;
			23427: outdata = 32'd42109;
			23428: outdata = 32'd42108;
			23429: outdata = 32'd42107;
			23430: outdata = 32'd42106;
			23431: outdata = 32'd42105;
			23432: outdata = 32'd42104;
			23433: outdata = 32'd42103;
			23434: outdata = 32'd42102;
			23435: outdata = 32'd42101;
			23436: outdata = 32'd42100;
			23437: outdata = 32'd42099;
			23438: outdata = 32'd42098;
			23439: outdata = 32'd42097;
			23440: outdata = 32'd42096;
			23441: outdata = 32'd42095;
			23442: outdata = 32'd42094;
			23443: outdata = 32'd42093;
			23444: outdata = 32'd42092;
			23445: outdata = 32'd42091;
			23446: outdata = 32'd42090;
			23447: outdata = 32'd42089;
			23448: outdata = 32'd42088;
			23449: outdata = 32'd42087;
			23450: outdata = 32'd42086;
			23451: outdata = 32'd42085;
			23452: outdata = 32'd42084;
			23453: outdata = 32'd42083;
			23454: outdata = 32'd42082;
			23455: outdata = 32'd42081;
			23456: outdata = 32'd42080;
			23457: outdata = 32'd42079;
			23458: outdata = 32'd42078;
			23459: outdata = 32'd42077;
			23460: outdata = 32'd42076;
			23461: outdata = 32'd42075;
			23462: outdata = 32'd42074;
			23463: outdata = 32'd42073;
			23464: outdata = 32'd42072;
			23465: outdata = 32'd42071;
			23466: outdata = 32'd42070;
			23467: outdata = 32'd42069;
			23468: outdata = 32'd42068;
			23469: outdata = 32'd42067;
			23470: outdata = 32'd42066;
			23471: outdata = 32'd42065;
			23472: outdata = 32'd42064;
			23473: outdata = 32'd42063;
			23474: outdata = 32'd42062;
			23475: outdata = 32'd42061;
			23476: outdata = 32'd42060;
			23477: outdata = 32'd42059;
			23478: outdata = 32'd42058;
			23479: outdata = 32'd42057;
			23480: outdata = 32'd42056;
			23481: outdata = 32'd42055;
			23482: outdata = 32'd42054;
			23483: outdata = 32'd42053;
			23484: outdata = 32'd42052;
			23485: outdata = 32'd42051;
			23486: outdata = 32'd42050;
			23487: outdata = 32'd42049;
			23488: outdata = 32'd42048;
			23489: outdata = 32'd42047;
			23490: outdata = 32'd42046;
			23491: outdata = 32'd42045;
			23492: outdata = 32'd42044;
			23493: outdata = 32'd42043;
			23494: outdata = 32'd42042;
			23495: outdata = 32'd42041;
			23496: outdata = 32'd42040;
			23497: outdata = 32'd42039;
			23498: outdata = 32'd42038;
			23499: outdata = 32'd42037;
			23500: outdata = 32'd42036;
			23501: outdata = 32'd42035;
			23502: outdata = 32'd42034;
			23503: outdata = 32'd42033;
			23504: outdata = 32'd42032;
			23505: outdata = 32'd42031;
			23506: outdata = 32'd42030;
			23507: outdata = 32'd42029;
			23508: outdata = 32'd42028;
			23509: outdata = 32'd42027;
			23510: outdata = 32'd42026;
			23511: outdata = 32'd42025;
			23512: outdata = 32'd42024;
			23513: outdata = 32'd42023;
			23514: outdata = 32'd42022;
			23515: outdata = 32'd42021;
			23516: outdata = 32'd42020;
			23517: outdata = 32'd42019;
			23518: outdata = 32'd42018;
			23519: outdata = 32'd42017;
			23520: outdata = 32'd42016;
			23521: outdata = 32'd42015;
			23522: outdata = 32'd42014;
			23523: outdata = 32'd42013;
			23524: outdata = 32'd42012;
			23525: outdata = 32'd42011;
			23526: outdata = 32'd42010;
			23527: outdata = 32'd42009;
			23528: outdata = 32'd42008;
			23529: outdata = 32'd42007;
			23530: outdata = 32'd42006;
			23531: outdata = 32'd42005;
			23532: outdata = 32'd42004;
			23533: outdata = 32'd42003;
			23534: outdata = 32'd42002;
			23535: outdata = 32'd42001;
			23536: outdata = 32'd42000;
			23537: outdata = 32'd41999;
			23538: outdata = 32'd41998;
			23539: outdata = 32'd41997;
			23540: outdata = 32'd41996;
			23541: outdata = 32'd41995;
			23542: outdata = 32'd41994;
			23543: outdata = 32'd41993;
			23544: outdata = 32'd41992;
			23545: outdata = 32'd41991;
			23546: outdata = 32'd41990;
			23547: outdata = 32'd41989;
			23548: outdata = 32'd41988;
			23549: outdata = 32'd41987;
			23550: outdata = 32'd41986;
			23551: outdata = 32'd41985;
			23552: outdata = 32'd41984;
			23553: outdata = 32'd41983;
			23554: outdata = 32'd41982;
			23555: outdata = 32'd41981;
			23556: outdata = 32'd41980;
			23557: outdata = 32'd41979;
			23558: outdata = 32'd41978;
			23559: outdata = 32'd41977;
			23560: outdata = 32'd41976;
			23561: outdata = 32'd41975;
			23562: outdata = 32'd41974;
			23563: outdata = 32'd41973;
			23564: outdata = 32'd41972;
			23565: outdata = 32'd41971;
			23566: outdata = 32'd41970;
			23567: outdata = 32'd41969;
			23568: outdata = 32'd41968;
			23569: outdata = 32'd41967;
			23570: outdata = 32'd41966;
			23571: outdata = 32'd41965;
			23572: outdata = 32'd41964;
			23573: outdata = 32'd41963;
			23574: outdata = 32'd41962;
			23575: outdata = 32'd41961;
			23576: outdata = 32'd41960;
			23577: outdata = 32'd41959;
			23578: outdata = 32'd41958;
			23579: outdata = 32'd41957;
			23580: outdata = 32'd41956;
			23581: outdata = 32'd41955;
			23582: outdata = 32'd41954;
			23583: outdata = 32'd41953;
			23584: outdata = 32'd41952;
			23585: outdata = 32'd41951;
			23586: outdata = 32'd41950;
			23587: outdata = 32'd41949;
			23588: outdata = 32'd41948;
			23589: outdata = 32'd41947;
			23590: outdata = 32'd41946;
			23591: outdata = 32'd41945;
			23592: outdata = 32'd41944;
			23593: outdata = 32'd41943;
			23594: outdata = 32'd41942;
			23595: outdata = 32'd41941;
			23596: outdata = 32'd41940;
			23597: outdata = 32'd41939;
			23598: outdata = 32'd41938;
			23599: outdata = 32'd41937;
			23600: outdata = 32'd41936;
			23601: outdata = 32'd41935;
			23602: outdata = 32'd41934;
			23603: outdata = 32'd41933;
			23604: outdata = 32'd41932;
			23605: outdata = 32'd41931;
			23606: outdata = 32'd41930;
			23607: outdata = 32'd41929;
			23608: outdata = 32'd41928;
			23609: outdata = 32'd41927;
			23610: outdata = 32'd41926;
			23611: outdata = 32'd41925;
			23612: outdata = 32'd41924;
			23613: outdata = 32'd41923;
			23614: outdata = 32'd41922;
			23615: outdata = 32'd41921;
			23616: outdata = 32'd41920;
			23617: outdata = 32'd41919;
			23618: outdata = 32'd41918;
			23619: outdata = 32'd41917;
			23620: outdata = 32'd41916;
			23621: outdata = 32'd41915;
			23622: outdata = 32'd41914;
			23623: outdata = 32'd41913;
			23624: outdata = 32'd41912;
			23625: outdata = 32'd41911;
			23626: outdata = 32'd41910;
			23627: outdata = 32'd41909;
			23628: outdata = 32'd41908;
			23629: outdata = 32'd41907;
			23630: outdata = 32'd41906;
			23631: outdata = 32'd41905;
			23632: outdata = 32'd41904;
			23633: outdata = 32'd41903;
			23634: outdata = 32'd41902;
			23635: outdata = 32'd41901;
			23636: outdata = 32'd41900;
			23637: outdata = 32'd41899;
			23638: outdata = 32'd41898;
			23639: outdata = 32'd41897;
			23640: outdata = 32'd41896;
			23641: outdata = 32'd41895;
			23642: outdata = 32'd41894;
			23643: outdata = 32'd41893;
			23644: outdata = 32'd41892;
			23645: outdata = 32'd41891;
			23646: outdata = 32'd41890;
			23647: outdata = 32'd41889;
			23648: outdata = 32'd41888;
			23649: outdata = 32'd41887;
			23650: outdata = 32'd41886;
			23651: outdata = 32'd41885;
			23652: outdata = 32'd41884;
			23653: outdata = 32'd41883;
			23654: outdata = 32'd41882;
			23655: outdata = 32'd41881;
			23656: outdata = 32'd41880;
			23657: outdata = 32'd41879;
			23658: outdata = 32'd41878;
			23659: outdata = 32'd41877;
			23660: outdata = 32'd41876;
			23661: outdata = 32'd41875;
			23662: outdata = 32'd41874;
			23663: outdata = 32'd41873;
			23664: outdata = 32'd41872;
			23665: outdata = 32'd41871;
			23666: outdata = 32'd41870;
			23667: outdata = 32'd41869;
			23668: outdata = 32'd41868;
			23669: outdata = 32'd41867;
			23670: outdata = 32'd41866;
			23671: outdata = 32'd41865;
			23672: outdata = 32'd41864;
			23673: outdata = 32'd41863;
			23674: outdata = 32'd41862;
			23675: outdata = 32'd41861;
			23676: outdata = 32'd41860;
			23677: outdata = 32'd41859;
			23678: outdata = 32'd41858;
			23679: outdata = 32'd41857;
			23680: outdata = 32'd41856;
			23681: outdata = 32'd41855;
			23682: outdata = 32'd41854;
			23683: outdata = 32'd41853;
			23684: outdata = 32'd41852;
			23685: outdata = 32'd41851;
			23686: outdata = 32'd41850;
			23687: outdata = 32'd41849;
			23688: outdata = 32'd41848;
			23689: outdata = 32'd41847;
			23690: outdata = 32'd41846;
			23691: outdata = 32'd41845;
			23692: outdata = 32'd41844;
			23693: outdata = 32'd41843;
			23694: outdata = 32'd41842;
			23695: outdata = 32'd41841;
			23696: outdata = 32'd41840;
			23697: outdata = 32'd41839;
			23698: outdata = 32'd41838;
			23699: outdata = 32'd41837;
			23700: outdata = 32'd41836;
			23701: outdata = 32'd41835;
			23702: outdata = 32'd41834;
			23703: outdata = 32'd41833;
			23704: outdata = 32'd41832;
			23705: outdata = 32'd41831;
			23706: outdata = 32'd41830;
			23707: outdata = 32'd41829;
			23708: outdata = 32'd41828;
			23709: outdata = 32'd41827;
			23710: outdata = 32'd41826;
			23711: outdata = 32'd41825;
			23712: outdata = 32'd41824;
			23713: outdata = 32'd41823;
			23714: outdata = 32'd41822;
			23715: outdata = 32'd41821;
			23716: outdata = 32'd41820;
			23717: outdata = 32'd41819;
			23718: outdata = 32'd41818;
			23719: outdata = 32'd41817;
			23720: outdata = 32'd41816;
			23721: outdata = 32'd41815;
			23722: outdata = 32'd41814;
			23723: outdata = 32'd41813;
			23724: outdata = 32'd41812;
			23725: outdata = 32'd41811;
			23726: outdata = 32'd41810;
			23727: outdata = 32'd41809;
			23728: outdata = 32'd41808;
			23729: outdata = 32'd41807;
			23730: outdata = 32'd41806;
			23731: outdata = 32'd41805;
			23732: outdata = 32'd41804;
			23733: outdata = 32'd41803;
			23734: outdata = 32'd41802;
			23735: outdata = 32'd41801;
			23736: outdata = 32'd41800;
			23737: outdata = 32'd41799;
			23738: outdata = 32'd41798;
			23739: outdata = 32'd41797;
			23740: outdata = 32'd41796;
			23741: outdata = 32'd41795;
			23742: outdata = 32'd41794;
			23743: outdata = 32'd41793;
			23744: outdata = 32'd41792;
			23745: outdata = 32'd41791;
			23746: outdata = 32'd41790;
			23747: outdata = 32'd41789;
			23748: outdata = 32'd41788;
			23749: outdata = 32'd41787;
			23750: outdata = 32'd41786;
			23751: outdata = 32'd41785;
			23752: outdata = 32'd41784;
			23753: outdata = 32'd41783;
			23754: outdata = 32'd41782;
			23755: outdata = 32'd41781;
			23756: outdata = 32'd41780;
			23757: outdata = 32'd41779;
			23758: outdata = 32'd41778;
			23759: outdata = 32'd41777;
			23760: outdata = 32'd41776;
			23761: outdata = 32'd41775;
			23762: outdata = 32'd41774;
			23763: outdata = 32'd41773;
			23764: outdata = 32'd41772;
			23765: outdata = 32'd41771;
			23766: outdata = 32'd41770;
			23767: outdata = 32'd41769;
			23768: outdata = 32'd41768;
			23769: outdata = 32'd41767;
			23770: outdata = 32'd41766;
			23771: outdata = 32'd41765;
			23772: outdata = 32'd41764;
			23773: outdata = 32'd41763;
			23774: outdata = 32'd41762;
			23775: outdata = 32'd41761;
			23776: outdata = 32'd41760;
			23777: outdata = 32'd41759;
			23778: outdata = 32'd41758;
			23779: outdata = 32'd41757;
			23780: outdata = 32'd41756;
			23781: outdata = 32'd41755;
			23782: outdata = 32'd41754;
			23783: outdata = 32'd41753;
			23784: outdata = 32'd41752;
			23785: outdata = 32'd41751;
			23786: outdata = 32'd41750;
			23787: outdata = 32'd41749;
			23788: outdata = 32'd41748;
			23789: outdata = 32'd41747;
			23790: outdata = 32'd41746;
			23791: outdata = 32'd41745;
			23792: outdata = 32'd41744;
			23793: outdata = 32'd41743;
			23794: outdata = 32'd41742;
			23795: outdata = 32'd41741;
			23796: outdata = 32'd41740;
			23797: outdata = 32'd41739;
			23798: outdata = 32'd41738;
			23799: outdata = 32'd41737;
			23800: outdata = 32'd41736;
			23801: outdata = 32'd41735;
			23802: outdata = 32'd41734;
			23803: outdata = 32'd41733;
			23804: outdata = 32'd41732;
			23805: outdata = 32'd41731;
			23806: outdata = 32'd41730;
			23807: outdata = 32'd41729;
			23808: outdata = 32'd41728;
			23809: outdata = 32'd41727;
			23810: outdata = 32'd41726;
			23811: outdata = 32'd41725;
			23812: outdata = 32'd41724;
			23813: outdata = 32'd41723;
			23814: outdata = 32'd41722;
			23815: outdata = 32'd41721;
			23816: outdata = 32'd41720;
			23817: outdata = 32'd41719;
			23818: outdata = 32'd41718;
			23819: outdata = 32'd41717;
			23820: outdata = 32'd41716;
			23821: outdata = 32'd41715;
			23822: outdata = 32'd41714;
			23823: outdata = 32'd41713;
			23824: outdata = 32'd41712;
			23825: outdata = 32'd41711;
			23826: outdata = 32'd41710;
			23827: outdata = 32'd41709;
			23828: outdata = 32'd41708;
			23829: outdata = 32'd41707;
			23830: outdata = 32'd41706;
			23831: outdata = 32'd41705;
			23832: outdata = 32'd41704;
			23833: outdata = 32'd41703;
			23834: outdata = 32'd41702;
			23835: outdata = 32'd41701;
			23836: outdata = 32'd41700;
			23837: outdata = 32'd41699;
			23838: outdata = 32'd41698;
			23839: outdata = 32'd41697;
			23840: outdata = 32'd41696;
			23841: outdata = 32'd41695;
			23842: outdata = 32'd41694;
			23843: outdata = 32'd41693;
			23844: outdata = 32'd41692;
			23845: outdata = 32'd41691;
			23846: outdata = 32'd41690;
			23847: outdata = 32'd41689;
			23848: outdata = 32'd41688;
			23849: outdata = 32'd41687;
			23850: outdata = 32'd41686;
			23851: outdata = 32'd41685;
			23852: outdata = 32'd41684;
			23853: outdata = 32'd41683;
			23854: outdata = 32'd41682;
			23855: outdata = 32'd41681;
			23856: outdata = 32'd41680;
			23857: outdata = 32'd41679;
			23858: outdata = 32'd41678;
			23859: outdata = 32'd41677;
			23860: outdata = 32'd41676;
			23861: outdata = 32'd41675;
			23862: outdata = 32'd41674;
			23863: outdata = 32'd41673;
			23864: outdata = 32'd41672;
			23865: outdata = 32'd41671;
			23866: outdata = 32'd41670;
			23867: outdata = 32'd41669;
			23868: outdata = 32'd41668;
			23869: outdata = 32'd41667;
			23870: outdata = 32'd41666;
			23871: outdata = 32'd41665;
			23872: outdata = 32'd41664;
			23873: outdata = 32'd41663;
			23874: outdata = 32'd41662;
			23875: outdata = 32'd41661;
			23876: outdata = 32'd41660;
			23877: outdata = 32'd41659;
			23878: outdata = 32'd41658;
			23879: outdata = 32'd41657;
			23880: outdata = 32'd41656;
			23881: outdata = 32'd41655;
			23882: outdata = 32'd41654;
			23883: outdata = 32'd41653;
			23884: outdata = 32'd41652;
			23885: outdata = 32'd41651;
			23886: outdata = 32'd41650;
			23887: outdata = 32'd41649;
			23888: outdata = 32'd41648;
			23889: outdata = 32'd41647;
			23890: outdata = 32'd41646;
			23891: outdata = 32'd41645;
			23892: outdata = 32'd41644;
			23893: outdata = 32'd41643;
			23894: outdata = 32'd41642;
			23895: outdata = 32'd41641;
			23896: outdata = 32'd41640;
			23897: outdata = 32'd41639;
			23898: outdata = 32'd41638;
			23899: outdata = 32'd41637;
			23900: outdata = 32'd41636;
			23901: outdata = 32'd41635;
			23902: outdata = 32'd41634;
			23903: outdata = 32'd41633;
			23904: outdata = 32'd41632;
			23905: outdata = 32'd41631;
			23906: outdata = 32'd41630;
			23907: outdata = 32'd41629;
			23908: outdata = 32'd41628;
			23909: outdata = 32'd41627;
			23910: outdata = 32'd41626;
			23911: outdata = 32'd41625;
			23912: outdata = 32'd41624;
			23913: outdata = 32'd41623;
			23914: outdata = 32'd41622;
			23915: outdata = 32'd41621;
			23916: outdata = 32'd41620;
			23917: outdata = 32'd41619;
			23918: outdata = 32'd41618;
			23919: outdata = 32'd41617;
			23920: outdata = 32'd41616;
			23921: outdata = 32'd41615;
			23922: outdata = 32'd41614;
			23923: outdata = 32'd41613;
			23924: outdata = 32'd41612;
			23925: outdata = 32'd41611;
			23926: outdata = 32'd41610;
			23927: outdata = 32'd41609;
			23928: outdata = 32'd41608;
			23929: outdata = 32'd41607;
			23930: outdata = 32'd41606;
			23931: outdata = 32'd41605;
			23932: outdata = 32'd41604;
			23933: outdata = 32'd41603;
			23934: outdata = 32'd41602;
			23935: outdata = 32'd41601;
			23936: outdata = 32'd41600;
			23937: outdata = 32'd41599;
			23938: outdata = 32'd41598;
			23939: outdata = 32'd41597;
			23940: outdata = 32'd41596;
			23941: outdata = 32'd41595;
			23942: outdata = 32'd41594;
			23943: outdata = 32'd41593;
			23944: outdata = 32'd41592;
			23945: outdata = 32'd41591;
			23946: outdata = 32'd41590;
			23947: outdata = 32'd41589;
			23948: outdata = 32'd41588;
			23949: outdata = 32'd41587;
			23950: outdata = 32'd41586;
			23951: outdata = 32'd41585;
			23952: outdata = 32'd41584;
			23953: outdata = 32'd41583;
			23954: outdata = 32'd41582;
			23955: outdata = 32'd41581;
			23956: outdata = 32'd41580;
			23957: outdata = 32'd41579;
			23958: outdata = 32'd41578;
			23959: outdata = 32'd41577;
			23960: outdata = 32'd41576;
			23961: outdata = 32'd41575;
			23962: outdata = 32'd41574;
			23963: outdata = 32'd41573;
			23964: outdata = 32'd41572;
			23965: outdata = 32'd41571;
			23966: outdata = 32'd41570;
			23967: outdata = 32'd41569;
			23968: outdata = 32'd41568;
			23969: outdata = 32'd41567;
			23970: outdata = 32'd41566;
			23971: outdata = 32'd41565;
			23972: outdata = 32'd41564;
			23973: outdata = 32'd41563;
			23974: outdata = 32'd41562;
			23975: outdata = 32'd41561;
			23976: outdata = 32'd41560;
			23977: outdata = 32'd41559;
			23978: outdata = 32'd41558;
			23979: outdata = 32'd41557;
			23980: outdata = 32'd41556;
			23981: outdata = 32'd41555;
			23982: outdata = 32'd41554;
			23983: outdata = 32'd41553;
			23984: outdata = 32'd41552;
			23985: outdata = 32'd41551;
			23986: outdata = 32'd41550;
			23987: outdata = 32'd41549;
			23988: outdata = 32'd41548;
			23989: outdata = 32'd41547;
			23990: outdata = 32'd41546;
			23991: outdata = 32'd41545;
			23992: outdata = 32'd41544;
			23993: outdata = 32'd41543;
			23994: outdata = 32'd41542;
			23995: outdata = 32'd41541;
			23996: outdata = 32'd41540;
			23997: outdata = 32'd41539;
			23998: outdata = 32'd41538;
			23999: outdata = 32'd41537;
			24000: outdata = 32'd41536;
			24001: outdata = 32'd41535;
			24002: outdata = 32'd41534;
			24003: outdata = 32'd41533;
			24004: outdata = 32'd41532;
			24005: outdata = 32'd41531;
			24006: outdata = 32'd41530;
			24007: outdata = 32'd41529;
			24008: outdata = 32'd41528;
			24009: outdata = 32'd41527;
			24010: outdata = 32'd41526;
			24011: outdata = 32'd41525;
			24012: outdata = 32'd41524;
			24013: outdata = 32'd41523;
			24014: outdata = 32'd41522;
			24015: outdata = 32'd41521;
			24016: outdata = 32'd41520;
			24017: outdata = 32'd41519;
			24018: outdata = 32'd41518;
			24019: outdata = 32'd41517;
			24020: outdata = 32'd41516;
			24021: outdata = 32'd41515;
			24022: outdata = 32'd41514;
			24023: outdata = 32'd41513;
			24024: outdata = 32'd41512;
			24025: outdata = 32'd41511;
			24026: outdata = 32'd41510;
			24027: outdata = 32'd41509;
			24028: outdata = 32'd41508;
			24029: outdata = 32'd41507;
			24030: outdata = 32'd41506;
			24031: outdata = 32'd41505;
			24032: outdata = 32'd41504;
			24033: outdata = 32'd41503;
			24034: outdata = 32'd41502;
			24035: outdata = 32'd41501;
			24036: outdata = 32'd41500;
			24037: outdata = 32'd41499;
			24038: outdata = 32'd41498;
			24039: outdata = 32'd41497;
			24040: outdata = 32'd41496;
			24041: outdata = 32'd41495;
			24042: outdata = 32'd41494;
			24043: outdata = 32'd41493;
			24044: outdata = 32'd41492;
			24045: outdata = 32'd41491;
			24046: outdata = 32'd41490;
			24047: outdata = 32'd41489;
			24048: outdata = 32'd41488;
			24049: outdata = 32'd41487;
			24050: outdata = 32'd41486;
			24051: outdata = 32'd41485;
			24052: outdata = 32'd41484;
			24053: outdata = 32'd41483;
			24054: outdata = 32'd41482;
			24055: outdata = 32'd41481;
			24056: outdata = 32'd41480;
			24057: outdata = 32'd41479;
			24058: outdata = 32'd41478;
			24059: outdata = 32'd41477;
			24060: outdata = 32'd41476;
			24061: outdata = 32'd41475;
			24062: outdata = 32'd41474;
			24063: outdata = 32'd41473;
			24064: outdata = 32'd41472;
			24065: outdata = 32'd41471;
			24066: outdata = 32'd41470;
			24067: outdata = 32'd41469;
			24068: outdata = 32'd41468;
			24069: outdata = 32'd41467;
			24070: outdata = 32'd41466;
			24071: outdata = 32'd41465;
			24072: outdata = 32'd41464;
			24073: outdata = 32'd41463;
			24074: outdata = 32'd41462;
			24075: outdata = 32'd41461;
			24076: outdata = 32'd41460;
			24077: outdata = 32'd41459;
			24078: outdata = 32'd41458;
			24079: outdata = 32'd41457;
			24080: outdata = 32'd41456;
			24081: outdata = 32'd41455;
			24082: outdata = 32'd41454;
			24083: outdata = 32'd41453;
			24084: outdata = 32'd41452;
			24085: outdata = 32'd41451;
			24086: outdata = 32'd41450;
			24087: outdata = 32'd41449;
			24088: outdata = 32'd41448;
			24089: outdata = 32'd41447;
			24090: outdata = 32'd41446;
			24091: outdata = 32'd41445;
			24092: outdata = 32'd41444;
			24093: outdata = 32'd41443;
			24094: outdata = 32'd41442;
			24095: outdata = 32'd41441;
			24096: outdata = 32'd41440;
			24097: outdata = 32'd41439;
			24098: outdata = 32'd41438;
			24099: outdata = 32'd41437;
			24100: outdata = 32'd41436;
			24101: outdata = 32'd41435;
			24102: outdata = 32'd41434;
			24103: outdata = 32'd41433;
			24104: outdata = 32'd41432;
			24105: outdata = 32'd41431;
			24106: outdata = 32'd41430;
			24107: outdata = 32'd41429;
			24108: outdata = 32'd41428;
			24109: outdata = 32'd41427;
			24110: outdata = 32'd41426;
			24111: outdata = 32'd41425;
			24112: outdata = 32'd41424;
			24113: outdata = 32'd41423;
			24114: outdata = 32'd41422;
			24115: outdata = 32'd41421;
			24116: outdata = 32'd41420;
			24117: outdata = 32'd41419;
			24118: outdata = 32'd41418;
			24119: outdata = 32'd41417;
			24120: outdata = 32'd41416;
			24121: outdata = 32'd41415;
			24122: outdata = 32'd41414;
			24123: outdata = 32'd41413;
			24124: outdata = 32'd41412;
			24125: outdata = 32'd41411;
			24126: outdata = 32'd41410;
			24127: outdata = 32'd41409;
			24128: outdata = 32'd41408;
			24129: outdata = 32'd41407;
			24130: outdata = 32'd41406;
			24131: outdata = 32'd41405;
			24132: outdata = 32'd41404;
			24133: outdata = 32'd41403;
			24134: outdata = 32'd41402;
			24135: outdata = 32'd41401;
			24136: outdata = 32'd41400;
			24137: outdata = 32'd41399;
			24138: outdata = 32'd41398;
			24139: outdata = 32'd41397;
			24140: outdata = 32'd41396;
			24141: outdata = 32'd41395;
			24142: outdata = 32'd41394;
			24143: outdata = 32'd41393;
			24144: outdata = 32'd41392;
			24145: outdata = 32'd41391;
			24146: outdata = 32'd41390;
			24147: outdata = 32'd41389;
			24148: outdata = 32'd41388;
			24149: outdata = 32'd41387;
			24150: outdata = 32'd41386;
			24151: outdata = 32'd41385;
			24152: outdata = 32'd41384;
			24153: outdata = 32'd41383;
			24154: outdata = 32'd41382;
			24155: outdata = 32'd41381;
			24156: outdata = 32'd41380;
			24157: outdata = 32'd41379;
			24158: outdata = 32'd41378;
			24159: outdata = 32'd41377;
			24160: outdata = 32'd41376;
			24161: outdata = 32'd41375;
			24162: outdata = 32'd41374;
			24163: outdata = 32'd41373;
			24164: outdata = 32'd41372;
			24165: outdata = 32'd41371;
			24166: outdata = 32'd41370;
			24167: outdata = 32'd41369;
			24168: outdata = 32'd41368;
			24169: outdata = 32'd41367;
			24170: outdata = 32'd41366;
			24171: outdata = 32'd41365;
			24172: outdata = 32'd41364;
			24173: outdata = 32'd41363;
			24174: outdata = 32'd41362;
			24175: outdata = 32'd41361;
			24176: outdata = 32'd41360;
			24177: outdata = 32'd41359;
			24178: outdata = 32'd41358;
			24179: outdata = 32'd41357;
			24180: outdata = 32'd41356;
			24181: outdata = 32'd41355;
			24182: outdata = 32'd41354;
			24183: outdata = 32'd41353;
			24184: outdata = 32'd41352;
			24185: outdata = 32'd41351;
			24186: outdata = 32'd41350;
			24187: outdata = 32'd41349;
			24188: outdata = 32'd41348;
			24189: outdata = 32'd41347;
			24190: outdata = 32'd41346;
			24191: outdata = 32'd41345;
			24192: outdata = 32'd41344;
			24193: outdata = 32'd41343;
			24194: outdata = 32'd41342;
			24195: outdata = 32'd41341;
			24196: outdata = 32'd41340;
			24197: outdata = 32'd41339;
			24198: outdata = 32'd41338;
			24199: outdata = 32'd41337;
			24200: outdata = 32'd41336;
			24201: outdata = 32'd41335;
			24202: outdata = 32'd41334;
			24203: outdata = 32'd41333;
			24204: outdata = 32'd41332;
			24205: outdata = 32'd41331;
			24206: outdata = 32'd41330;
			24207: outdata = 32'd41329;
			24208: outdata = 32'd41328;
			24209: outdata = 32'd41327;
			24210: outdata = 32'd41326;
			24211: outdata = 32'd41325;
			24212: outdata = 32'd41324;
			24213: outdata = 32'd41323;
			24214: outdata = 32'd41322;
			24215: outdata = 32'd41321;
			24216: outdata = 32'd41320;
			24217: outdata = 32'd41319;
			24218: outdata = 32'd41318;
			24219: outdata = 32'd41317;
			24220: outdata = 32'd41316;
			24221: outdata = 32'd41315;
			24222: outdata = 32'd41314;
			24223: outdata = 32'd41313;
			24224: outdata = 32'd41312;
			24225: outdata = 32'd41311;
			24226: outdata = 32'd41310;
			24227: outdata = 32'd41309;
			24228: outdata = 32'd41308;
			24229: outdata = 32'd41307;
			24230: outdata = 32'd41306;
			24231: outdata = 32'd41305;
			24232: outdata = 32'd41304;
			24233: outdata = 32'd41303;
			24234: outdata = 32'd41302;
			24235: outdata = 32'd41301;
			24236: outdata = 32'd41300;
			24237: outdata = 32'd41299;
			24238: outdata = 32'd41298;
			24239: outdata = 32'd41297;
			24240: outdata = 32'd41296;
			24241: outdata = 32'd41295;
			24242: outdata = 32'd41294;
			24243: outdata = 32'd41293;
			24244: outdata = 32'd41292;
			24245: outdata = 32'd41291;
			24246: outdata = 32'd41290;
			24247: outdata = 32'd41289;
			24248: outdata = 32'd41288;
			24249: outdata = 32'd41287;
			24250: outdata = 32'd41286;
			24251: outdata = 32'd41285;
			24252: outdata = 32'd41284;
			24253: outdata = 32'd41283;
			24254: outdata = 32'd41282;
			24255: outdata = 32'd41281;
			24256: outdata = 32'd41280;
			24257: outdata = 32'd41279;
			24258: outdata = 32'd41278;
			24259: outdata = 32'd41277;
			24260: outdata = 32'd41276;
			24261: outdata = 32'd41275;
			24262: outdata = 32'd41274;
			24263: outdata = 32'd41273;
			24264: outdata = 32'd41272;
			24265: outdata = 32'd41271;
			24266: outdata = 32'd41270;
			24267: outdata = 32'd41269;
			24268: outdata = 32'd41268;
			24269: outdata = 32'd41267;
			24270: outdata = 32'd41266;
			24271: outdata = 32'd41265;
			24272: outdata = 32'd41264;
			24273: outdata = 32'd41263;
			24274: outdata = 32'd41262;
			24275: outdata = 32'd41261;
			24276: outdata = 32'd41260;
			24277: outdata = 32'd41259;
			24278: outdata = 32'd41258;
			24279: outdata = 32'd41257;
			24280: outdata = 32'd41256;
			24281: outdata = 32'd41255;
			24282: outdata = 32'd41254;
			24283: outdata = 32'd41253;
			24284: outdata = 32'd41252;
			24285: outdata = 32'd41251;
			24286: outdata = 32'd41250;
			24287: outdata = 32'd41249;
			24288: outdata = 32'd41248;
			24289: outdata = 32'd41247;
			24290: outdata = 32'd41246;
			24291: outdata = 32'd41245;
			24292: outdata = 32'd41244;
			24293: outdata = 32'd41243;
			24294: outdata = 32'd41242;
			24295: outdata = 32'd41241;
			24296: outdata = 32'd41240;
			24297: outdata = 32'd41239;
			24298: outdata = 32'd41238;
			24299: outdata = 32'd41237;
			24300: outdata = 32'd41236;
			24301: outdata = 32'd41235;
			24302: outdata = 32'd41234;
			24303: outdata = 32'd41233;
			24304: outdata = 32'd41232;
			24305: outdata = 32'd41231;
			24306: outdata = 32'd41230;
			24307: outdata = 32'd41229;
			24308: outdata = 32'd41228;
			24309: outdata = 32'd41227;
			24310: outdata = 32'd41226;
			24311: outdata = 32'd41225;
			24312: outdata = 32'd41224;
			24313: outdata = 32'd41223;
			24314: outdata = 32'd41222;
			24315: outdata = 32'd41221;
			24316: outdata = 32'd41220;
			24317: outdata = 32'd41219;
			24318: outdata = 32'd41218;
			24319: outdata = 32'd41217;
			24320: outdata = 32'd41216;
			24321: outdata = 32'd41215;
			24322: outdata = 32'd41214;
			24323: outdata = 32'd41213;
			24324: outdata = 32'd41212;
			24325: outdata = 32'd41211;
			24326: outdata = 32'd41210;
			24327: outdata = 32'd41209;
			24328: outdata = 32'd41208;
			24329: outdata = 32'd41207;
			24330: outdata = 32'd41206;
			24331: outdata = 32'd41205;
			24332: outdata = 32'd41204;
			24333: outdata = 32'd41203;
			24334: outdata = 32'd41202;
			24335: outdata = 32'd41201;
			24336: outdata = 32'd41200;
			24337: outdata = 32'd41199;
			24338: outdata = 32'd41198;
			24339: outdata = 32'd41197;
			24340: outdata = 32'd41196;
			24341: outdata = 32'd41195;
			24342: outdata = 32'd41194;
			24343: outdata = 32'd41193;
			24344: outdata = 32'd41192;
			24345: outdata = 32'd41191;
			24346: outdata = 32'd41190;
			24347: outdata = 32'd41189;
			24348: outdata = 32'd41188;
			24349: outdata = 32'd41187;
			24350: outdata = 32'd41186;
			24351: outdata = 32'd41185;
			24352: outdata = 32'd41184;
			24353: outdata = 32'd41183;
			24354: outdata = 32'd41182;
			24355: outdata = 32'd41181;
			24356: outdata = 32'd41180;
			24357: outdata = 32'd41179;
			24358: outdata = 32'd41178;
			24359: outdata = 32'd41177;
			24360: outdata = 32'd41176;
			24361: outdata = 32'd41175;
			24362: outdata = 32'd41174;
			24363: outdata = 32'd41173;
			24364: outdata = 32'd41172;
			24365: outdata = 32'd41171;
			24366: outdata = 32'd41170;
			24367: outdata = 32'd41169;
			24368: outdata = 32'd41168;
			24369: outdata = 32'd41167;
			24370: outdata = 32'd41166;
			24371: outdata = 32'd41165;
			24372: outdata = 32'd41164;
			24373: outdata = 32'd41163;
			24374: outdata = 32'd41162;
			24375: outdata = 32'd41161;
			24376: outdata = 32'd41160;
			24377: outdata = 32'd41159;
			24378: outdata = 32'd41158;
			24379: outdata = 32'd41157;
			24380: outdata = 32'd41156;
			24381: outdata = 32'd41155;
			24382: outdata = 32'd41154;
			24383: outdata = 32'd41153;
			24384: outdata = 32'd41152;
			24385: outdata = 32'd41151;
			24386: outdata = 32'd41150;
			24387: outdata = 32'd41149;
			24388: outdata = 32'd41148;
			24389: outdata = 32'd41147;
			24390: outdata = 32'd41146;
			24391: outdata = 32'd41145;
			24392: outdata = 32'd41144;
			24393: outdata = 32'd41143;
			24394: outdata = 32'd41142;
			24395: outdata = 32'd41141;
			24396: outdata = 32'd41140;
			24397: outdata = 32'd41139;
			24398: outdata = 32'd41138;
			24399: outdata = 32'd41137;
			24400: outdata = 32'd41136;
			24401: outdata = 32'd41135;
			24402: outdata = 32'd41134;
			24403: outdata = 32'd41133;
			24404: outdata = 32'd41132;
			24405: outdata = 32'd41131;
			24406: outdata = 32'd41130;
			24407: outdata = 32'd41129;
			24408: outdata = 32'd41128;
			24409: outdata = 32'd41127;
			24410: outdata = 32'd41126;
			24411: outdata = 32'd41125;
			24412: outdata = 32'd41124;
			24413: outdata = 32'd41123;
			24414: outdata = 32'd41122;
			24415: outdata = 32'd41121;
			24416: outdata = 32'd41120;
			24417: outdata = 32'd41119;
			24418: outdata = 32'd41118;
			24419: outdata = 32'd41117;
			24420: outdata = 32'd41116;
			24421: outdata = 32'd41115;
			24422: outdata = 32'd41114;
			24423: outdata = 32'd41113;
			24424: outdata = 32'd41112;
			24425: outdata = 32'd41111;
			24426: outdata = 32'd41110;
			24427: outdata = 32'd41109;
			24428: outdata = 32'd41108;
			24429: outdata = 32'd41107;
			24430: outdata = 32'd41106;
			24431: outdata = 32'd41105;
			24432: outdata = 32'd41104;
			24433: outdata = 32'd41103;
			24434: outdata = 32'd41102;
			24435: outdata = 32'd41101;
			24436: outdata = 32'd41100;
			24437: outdata = 32'd41099;
			24438: outdata = 32'd41098;
			24439: outdata = 32'd41097;
			24440: outdata = 32'd41096;
			24441: outdata = 32'd41095;
			24442: outdata = 32'd41094;
			24443: outdata = 32'd41093;
			24444: outdata = 32'd41092;
			24445: outdata = 32'd41091;
			24446: outdata = 32'd41090;
			24447: outdata = 32'd41089;
			24448: outdata = 32'd41088;
			24449: outdata = 32'd41087;
			24450: outdata = 32'd41086;
			24451: outdata = 32'd41085;
			24452: outdata = 32'd41084;
			24453: outdata = 32'd41083;
			24454: outdata = 32'd41082;
			24455: outdata = 32'd41081;
			24456: outdata = 32'd41080;
			24457: outdata = 32'd41079;
			24458: outdata = 32'd41078;
			24459: outdata = 32'd41077;
			24460: outdata = 32'd41076;
			24461: outdata = 32'd41075;
			24462: outdata = 32'd41074;
			24463: outdata = 32'd41073;
			24464: outdata = 32'd41072;
			24465: outdata = 32'd41071;
			24466: outdata = 32'd41070;
			24467: outdata = 32'd41069;
			24468: outdata = 32'd41068;
			24469: outdata = 32'd41067;
			24470: outdata = 32'd41066;
			24471: outdata = 32'd41065;
			24472: outdata = 32'd41064;
			24473: outdata = 32'd41063;
			24474: outdata = 32'd41062;
			24475: outdata = 32'd41061;
			24476: outdata = 32'd41060;
			24477: outdata = 32'd41059;
			24478: outdata = 32'd41058;
			24479: outdata = 32'd41057;
			24480: outdata = 32'd41056;
			24481: outdata = 32'd41055;
			24482: outdata = 32'd41054;
			24483: outdata = 32'd41053;
			24484: outdata = 32'd41052;
			24485: outdata = 32'd41051;
			24486: outdata = 32'd41050;
			24487: outdata = 32'd41049;
			24488: outdata = 32'd41048;
			24489: outdata = 32'd41047;
			24490: outdata = 32'd41046;
			24491: outdata = 32'd41045;
			24492: outdata = 32'd41044;
			24493: outdata = 32'd41043;
			24494: outdata = 32'd41042;
			24495: outdata = 32'd41041;
			24496: outdata = 32'd41040;
			24497: outdata = 32'd41039;
			24498: outdata = 32'd41038;
			24499: outdata = 32'd41037;
			24500: outdata = 32'd41036;
			24501: outdata = 32'd41035;
			24502: outdata = 32'd41034;
			24503: outdata = 32'd41033;
			24504: outdata = 32'd41032;
			24505: outdata = 32'd41031;
			24506: outdata = 32'd41030;
			24507: outdata = 32'd41029;
			24508: outdata = 32'd41028;
			24509: outdata = 32'd41027;
			24510: outdata = 32'd41026;
			24511: outdata = 32'd41025;
			24512: outdata = 32'd41024;
			24513: outdata = 32'd41023;
			24514: outdata = 32'd41022;
			24515: outdata = 32'd41021;
			24516: outdata = 32'd41020;
			24517: outdata = 32'd41019;
			24518: outdata = 32'd41018;
			24519: outdata = 32'd41017;
			24520: outdata = 32'd41016;
			24521: outdata = 32'd41015;
			24522: outdata = 32'd41014;
			24523: outdata = 32'd41013;
			24524: outdata = 32'd41012;
			24525: outdata = 32'd41011;
			24526: outdata = 32'd41010;
			24527: outdata = 32'd41009;
			24528: outdata = 32'd41008;
			24529: outdata = 32'd41007;
			24530: outdata = 32'd41006;
			24531: outdata = 32'd41005;
			24532: outdata = 32'd41004;
			24533: outdata = 32'd41003;
			24534: outdata = 32'd41002;
			24535: outdata = 32'd41001;
			24536: outdata = 32'd41000;
			24537: outdata = 32'd40999;
			24538: outdata = 32'd40998;
			24539: outdata = 32'd40997;
			24540: outdata = 32'd40996;
			24541: outdata = 32'd40995;
			24542: outdata = 32'd40994;
			24543: outdata = 32'd40993;
			24544: outdata = 32'd40992;
			24545: outdata = 32'd40991;
			24546: outdata = 32'd40990;
			24547: outdata = 32'd40989;
			24548: outdata = 32'd40988;
			24549: outdata = 32'd40987;
			24550: outdata = 32'd40986;
			24551: outdata = 32'd40985;
			24552: outdata = 32'd40984;
			24553: outdata = 32'd40983;
			24554: outdata = 32'd40982;
			24555: outdata = 32'd40981;
			24556: outdata = 32'd40980;
			24557: outdata = 32'd40979;
			24558: outdata = 32'd40978;
			24559: outdata = 32'd40977;
			24560: outdata = 32'd40976;
			24561: outdata = 32'd40975;
			24562: outdata = 32'd40974;
			24563: outdata = 32'd40973;
			24564: outdata = 32'd40972;
			24565: outdata = 32'd40971;
			24566: outdata = 32'd40970;
			24567: outdata = 32'd40969;
			24568: outdata = 32'd40968;
			24569: outdata = 32'd40967;
			24570: outdata = 32'd40966;
			24571: outdata = 32'd40965;
			24572: outdata = 32'd40964;
			24573: outdata = 32'd40963;
			24574: outdata = 32'd40962;
			24575: outdata = 32'd40961;
			24576: outdata = 32'd40960;
			24577: outdata = 32'd40959;
			24578: outdata = 32'd40958;
			24579: outdata = 32'd40957;
			24580: outdata = 32'd40956;
			24581: outdata = 32'd40955;
			24582: outdata = 32'd40954;
			24583: outdata = 32'd40953;
			24584: outdata = 32'd40952;
			24585: outdata = 32'd40951;
			24586: outdata = 32'd40950;
			24587: outdata = 32'd40949;
			24588: outdata = 32'd40948;
			24589: outdata = 32'd40947;
			24590: outdata = 32'd40946;
			24591: outdata = 32'd40945;
			24592: outdata = 32'd40944;
			24593: outdata = 32'd40943;
			24594: outdata = 32'd40942;
			24595: outdata = 32'd40941;
			24596: outdata = 32'd40940;
			24597: outdata = 32'd40939;
			24598: outdata = 32'd40938;
			24599: outdata = 32'd40937;
			24600: outdata = 32'd40936;
			24601: outdata = 32'd40935;
			24602: outdata = 32'd40934;
			24603: outdata = 32'd40933;
			24604: outdata = 32'd40932;
			24605: outdata = 32'd40931;
			24606: outdata = 32'd40930;
			24607: outdata = 32'd40929;
			24608: outdata = 32'd40928;
			24609: outdata = 32'd40927;
			24610: outdata = 32'd40926;
			24611: outdata = 32'd40925;
			24612: outdata = 32'd40924;
			24613: outdata = 32'd40923;
			24614: outdata = 32'd40922;
			24615: outdata = 32'd40921;
			24616: outdata = 32'd40920;
			24617: outdata = 32'd40919;
			24618: outdata = 32'd40918;
			24619: outdata = 32'd40917;
			24620: outdata = 32'd40916;
			24621: outdata = 32'd40915;
			24622: outdata = 32'd40914;
			24623: outdata = 32'd40913;
			24624: outdata = 32'd40912;
			24625: outdata = 32'd40911;
			24626: outdata = 32'd40910;
			24627: outdata = 32'd40909;
			24628: outdata = 32'd40908;
			24629: outdata = 32'd40907;
			24630: outdata = 32'd40906;
			24631: outdata = 32'd40905;
			24632: outdata = 32'd40904;
			24633: outdata = 32'd40903;
			24634: outdata = 32'd40902;
			24635: outdata = 32'd40901;
			24636: outdata = 32'd40900;
			24637: outdata = 32'd40899;
			24638: outdata = 32'd40898;
			24639: outdata = 32'd40897;
			24640: outdata = 32'd40896;
			24641: outdata = 32'd40895;
			24642: outdata = 32'd40894;
			24643: outdata = 32'd40893;
			24644: outdata = 32'd40892;
			24645: outdata = 32'd40891;
			24646: outdata = 32'd40890;
			24647: outdata = 32'd40889;
			24648: outdata = 32'd40888;
			24649: outdata = 32'd40887;
			24650: outdata = 32'd40886;
			24651: outdata = 32'd40885;
			24652: outdata = 32'd40884;
			24653: outdata = 32'd40883;
			24654: outdata = 32'd40882;
			24655: outdata = 32'd40881;
			24656: outdata = 32'd40880;
			24657: outdata = 32'd40879;
			24658: outdata = 32'd40878;
			24659: outdata = 32'd40877;
			24660: outdata = 32'd40876;
			24661: outdata = 32'd40875;
			24662: outdata = 32'd40874;
			24663: outdata = 32'd40873;
			24664: outdata = 32'd40872;
			24665: outdata = 32'd40871;
			24666: outdata = 32'd40870;
			24667: outdata = 32'd40869;
			24668: outdata = 32'd40868;
			24669: outdata = 32'd40867;
			24670: outdata = 32'd40866;
			24671: outdata = 32'd40865;
			24672: outdata = 32'd40864;
			24673: outdata = 32'd40863;
			24674: outdata = 32'd40862;
			24675: outdata = 32'd40861;
			24676: outdata = 32'd40860;
			24677: outdata = 32'd40859;
			24678: outdata = 32'd40858;
			24679: outdata = 32'd40857;
			24680: outdata = 32'd40856;
			24681: outdata = 32'd40855;
			24682: outdata = 32'd40854;
			24683: outdata = 32'd40853;
			24684: outdata = 32'd40852;
			24685: outdata = 32'd40851;
			24686: outdata = 32'd40850;
			24687: outdata = 32'd40849;
			24688: outdata = 32'd40848;
			24689: outdata = 32'd40847;
			24690: outdata = 32'd40846;
			24691: outdata = 32'd40845;
			24692: outdata = 32'd40844;
			24693: outdata = 32'd40843;
			24694: outdata = 32'd40842;
			24695: outdata = 32'd40841;
			24696: outdata = 32'd40840;
			24697: outdata = 32'd40839;
			24698: outdata = 32'd40838;
			24699: outdata = 32'd40837;
			24700: outdata = 32'd40836;
			24701: outdata = 32'd40835;
			24702: outdata = 32'd40834;
			24703: outdata = 32'd40833;
			24704: outdata = 32'd40832;
			24705: outdata = 32'd40831;
			24706: outdata = 32'd40830;
			24707: outdata = 32'd40829;
			24708: outdata = 32'd40828;
			24709: outdata = 32'd40827;
			24710: outdata = 32'd40826;
			24711: outdata = 32'd40825;
			24712: outdata = 32'd40824;
			24713: outdata = 32'd40823;
			24714: outdata = 32'd40822;
			24715: outdata = 32'd40821;
			24716: outdata = 32'd40820;
			24717: outdata = 32'd40819;
			24718: outdata = 32'd40818;
			24719: outdata = 32'd40817;
			24720: outdata = 32'd40816;
			24721: outdata = 32'd40815;
			24722: outdata = 32'd40814;
			24723: outdata = 32'd40813;
			24724: outdata = 32'd40812;
			24725: outdata = 32'd40811;
			24726: outdata = 32'd40810;
			24727: outdata = 32'd40809;
			24728: outdata = 32'd40808;
			24729: outdata = 32'd40807;
			24730: outdata = 32'd40806;
			24731: outdata = 32'd40805;
			24732: outdata = 32'd40804;
			24733: outdata = 32'd40803;
			24734: outdata = 32'd40802;
			24735: outdata = 32'd40801;
			24736: outdata = 32'd40800;
			24737: outdata = 32'd40799;
			24738: outdata = 32'd40798;
			24739: outdata = 32'd40797;
			24740: outdata = 32'd40796;
			24741: outdata = 32'd40795;
			24742: outdata = 32'd40794;
			24743: outdata = 32'd40793;
			24744: outdata = 32'd40792;
			24745: outdata = 32'd40791;
			24746: outdata = 32'd40790;
			24747: outdata = 32'd40789;
			24748: outdata = 32'd40788;
			24749: outdata = 32'd40787;
			24750: outdata = 32'd40786;
			24751: outdata = 32'd40785;
			24752: outdata = 32'd40784;
			24753: outdata = 32'd40783;
			24754: outdata = 32'd40782;
			24755: outdata = 32'd40781;
			24756: outdata = 32'd40780;
			24757: outdata = 32'd40779;
			24758: outdata = 32'd40778;
			24759: outdata = 32'd40777;
			24760: outdata = 32'd40776;
			24761: outdata = 32'd40775;
			24762: outdata = 32'd40774;
			24763: outdata = 32'd40773;
			24764: outdata = 32'd40772;
			24765: outdata = 32'd40771;
			24766: outdata = 32'd40770;
			24767: outdata = 32'd40769;
			24768: outdata = 32'd40768;
			24769: outdata = 32'd40767;
			24770: outdata = 32'd40766;
			24771: outdata = 32'd40765;
			24772: outdata = 32'd40764;
			24773: outdata = 32'd40763;
			24774: outdata = 32'd40762;
			24775: outdata = 32'd40761;
			24776: outdata = 32'd40760;
			24777: outdata = 32'd40759;
			24778: outdata = 32'd40758;
			24779: outdata = 32'd40757;
			24780: outdata = 32'd40756;
			24781: outdata = 32'd40755;
			24782: outdata = 32'd40754;
			24783: outdata = 32'd40753;
			24784: outdata = 32'd40752;
			24785: outdata = 32'd40751;
			24786: outdata = 32'd40750;
			24787: outdata = 32'd40749;
			24788: outdata = 32'd40748;
			24789: outdata = 32'd40747;
			24790: outdata = 32'd40746;
			24791: outdata = 32'd40745;
			24792: outdata = 32'd40744;
			24793: outdata = 32'd40743;
			24794: outdata = 32'd40742;
			24795: outdata = 32'd40741;
			24796: outdata = 32'd40740;
			24797: outdata = 32'd40739;
			24798: outdata = 32'd40738;
			24799: outdata = 32'd40737;
			24800: outdata = 32'd40736;
			24801: outdata = 32'd40735;
			24802: outdata = 32'd40734;
			24803: outdata = 32'd40733;
			24804: outdata = 32'd40732;
			24805: outdata = 32'd40731;
			24806: outdata = 32'd40730;
			24807: outdata = 32'd40729;
			24808: outdata = 32'd40728;
			24809: outdata = 32'd40727;
			24810: outdata = 32'd40726;
			24811: outdata = 32'd40725;
			24812: outdata = 32'd40724;
			24813: outdata = 32'd40723;
			24814: outdata = 32'd40722;
			24815: outdata = 32'd40721;
			24816: outdata = 32'd40720;
			24817: outdata = 32'd40719;
			24818: outdata = 32'd40718;
			24819: outdata = 32'd40717;
			24820: outdata = 32'd40716;
			24821: outdata = 32'd40715;
			24822: outdata = 32'd40714;
			24823: outdata = 32'd40713;
			24824: outdata = 32'd40712;
			24825: outdata = 32'd40711;
			24826: outdata = 32'd40710;
			24827: outdata = 32'd40709;
			24828: outdata = 32'd40708;
			24829: outdata = 32'd40707;
			24830: outdata = 32'd40706;
			24831: outdata = 32'd40705;
			24832: outdata = 32'd40704;
			24833: outdata = 32'd40703;
			24834: outdata = 32'd40702;
			24835: outdata = 32'd40701;
			24836: outdata = 32'd40700;
			24837: outdata = 32'd40699;
			24838: outdata = 32'd40698;
			24839: outdata = 32'd40697;
			24840: outdata = 32'd40696;
			24841: outdata = 32'd40695;
			24842: outdata = 32'd40694;
			24843: outdata = 32'd40693;
			24844: outdata = 32'd40692;
			24845: outdata = 32'd40691;
			24846: outdata = 32'd40690;
			24847: outdata = 32'd40689;
			24848: outdata = 32'd40688;
			24849: outdata = 32'd40687;
			24850: outdata = 32'd40686;
			24851: outdata = 32'd40685;
			24852: outdata = 32'd40684;
			24853: outdata = 32'd40683;
			24854: outdata = 32'd40682;
			24855: outdata = 32'd40681;
			24856: outdata = 32'd40680;
			24857: outdata = 32'd40679;
			24858: outdata = 32'd40678;
			24859: outdata = 32'd40677;
			24860: outdata = 32'd40676;
			24861: outdata = 32'd40675;
			24862: outdata = 32'd40674;
			24863: outdata = 32'd40673;
			24864: outdata = 32'd40672;
			24865: outdata = 32'd40671;
			24866: outdata = 32'd40670;
			24867: outdata = 32'd40669;
			24868: outdata = 32'd40668;
			24869: outdata = 32'd40667;
			24870: outdata = 32'd40666;
			24871: outdata = 32'd40665;
			24872: outdata = 32'd40664;
			24873: outdata = 32'd40663;
			24874: outdata = 32'd40662;
			24875: outdata = 32'd40661;
			24876: outdata = 32'd40660;
			24877: outdata = 32'd40659;
			24878: outdata = 32'd40658;
			24879: outdata = 32'd40657;
			24880: outdata = 32'd40656;
			24881: outdata = 32'd40655;
			24882: outdata = 32'd40654;
			24883: outdata = 32'd40653;
			24884: outdata = 32'd40652;
			24885: outdata = 32'd40651;
			24886: outdata = 32'd40650;
			24887: outdata = 32'd40649;
			24888: outdata = 32'd40648;
			24889: outdata = 32'd40647;
			24890: outdata = 32'd40646;
			24891: outdata = 32'd40645;
			24892: outdata = 32'd40644;
			24893: outdata = 32'd40643;
			24894: outdata = 32'd40642;
			24895: outdata = 32'd40641;
			24896: outdata = 32'd40640;
			24897: outdata = 32'd40639;
			24898: outdata = 32'd40638;
			24899: outdata = 32'd40637;
			24900: outdata = 32'd40636;
			24901: outdata = 32'd40635;
			24902: outdata = 32'd40634;
			24903: outdata = 32'd40633;
			24904: outdata = 32'd40632;
			24905: outdata = 32'd40631;
			24906: outdata = 32'd40630;
			24907: outdata = 32'd40629;
			24908: outdata = 32'd40628;
			24909: outdata = 32'd40627;
			24910: outdata = 32'd40626;
			24911: outdata = 32'd40625;
			24912: outdata = 32'd40624;
			24913: outdata = 32'd40623;
			24914: outdata = 32'd40622;
			24915: outdata = 32'd40621;
			24916: outdata = 32'd40620;
			24917: outdata = 32'd40619;
			24918: outdata = 32'd40618;
			24919: outdata = 32'd40617;
			24920: outdata = 32'd40616;
			24921: outdata = 32'd40615;
			24922: outdata = 32'd40614;
			24923: outdata = 32'd40613;
			24924: outdata = 32'd40612;
			24925: outdata = 32'd40611;
			24926: outdata = 32'd40610;
			24927: outdata = 32'd40609;
			24928: outdata = 32'd40608;
			24929: outdata = 32'd40607;
			24930: outdata = 32'd40606;
			24931: outdata = 32'd40605;
			24932: outdata = 32'd40604;
			24933: outdata = 32'd40603;
			24934: outdata = 32'd40602;
			24935: outdata = 32'd40601;
			24936: outdata = 32'd40600;
			24937: outdata = 32'd40599;
			24938: outdata = 32'd40598;
			24939: outdata = 32'd40597;
			24940: outdata = 32'd40596;
			24941: outdata = 32'd40595;
			24942: outdata = 32'd40594;
			24943: outdata = 32'd40593;
			24944: outdata = 32'd40592;
			24945: outdata = 32'd40591;
			24946: outdata = 32'd40590;
			24947: outdata = 32'd40589;
			24948: outdata = 32'd40588;
			24949: outdata = 32'd40587;
			24950: outdata = 32'd40586;
			24951: outdata = 32'd40585;
			24952: outdata = 32'd40584;
			24953: outdata = 32'd40583;
			24954: outdata = 32'd40582;
			24955: outdata = 32'd40581;
			24956: outdata = 32'd40580;
			24957: outdata = 32'd40579;
			24958: outdata = 32'd40578;
			24959: outdata = 32'd40577;
			24960: outdata = 32'd40576;
			24961: outdata = 32'd40575;
			24962: outdata = 32'd40574;
			24963: outdata = 32'd40573;
			24964: outdata = 32'd40572;
			24965: outdata = 32'd40571;
			24966: outdata = 32'd40570;
			24967: outdata = 32'd40569;
			24968: outdata = 32'd40568;
			24969: outdata = 32'd40567;
			24970: outdata = 32'd40566;
			24971: outdata = 32'd40565;
			24972: outdata = 32'd40564;
			24973: outdata = 32'd40563;
			24974: outdata = 32'd40562;
			24975: outdata = 32'd40561;
			24976: outdata = 32'd40560;
			24977: outdata = 32'd40559;
			24978: outdata = 32'd40558;
			24979: outdata = 32'd40557;
			24980: outdata = 32'd40556;
			24981: outdata = 32'd40555;
			24982: outdata = 32'd40554;
			24983: outdata = 32'd40553;
			24984: outdata = 32'd40552;
			24985: outdata = 32'd40551;
			24986: outdata = 32'd40550;
			24987: outdata = 32'd40549;
			24988: outdata = 32'd40548;
			24989: outdata = 32'd40547;
			24990: outdata = 32'd40546;
			24991: outdata = 32'd40545;
			24992: outdata = 32'd40544;
			24993: outdata = 32'd40543;
			24994: outdata = 32'd40542;
			24995: outdata = 32'd40541;
			24996: outdata = 32'd40540;
			24997: outdata = 32'd40539;
			24998: outdata = 32'd40538;
			24999: outdata = 32'd40537;
			25000: outdata = 32'd40536;
			25001: outdata = 32'd40535;
			25002: outdata = 32'd40534;
			25003: outdata = 32'd40533;
			25004: outdata = 32'd40532;
			25005: outdata = 32'd40531;
			25006: outdata = 32'd40530;
			25007: outdata = 32'd40529;
			25008: outdata = 32'd40528;
			25009: outdata = 32'd40527;
			25010: outdata = 32'd40526;
			25011: outdata = 32'd40525;
			25012: outdata = 32'd40524;
			25013: outdata = 32'd40523;
			25014: outdata = 32'd40522;
			25015: outdata = 32'd40521;
			25016: outdata = 32'd40520;
			25017: outdata = 32'd40519;
			25018: outdata = 32'd40518;
			25019: outdata = 32'd40517;
			25020: outdata = 32'd40516;
			25021: outdata = 32'd40515;
			25022: outdata = 32'd40514;
			25023: outdata = 32'd40513;
			25024: outdata = 32'd40512;
			25025: outdata = 32'd40511;
			25026: outdata = 32'd40510;
			25027: outdata = 32'd40509;
			25028: outdata = 32'd40508;
			25029: outdata = 32'd40507;
			25030: outdata = 32'd40506;
			25031: outdata = 32'd40505;
			25032: outdata = 32'd40504;
			25033: outdata = 32'd40503;
			25034: outdata = 32'd40502;
			25035: outdata = 32'd40501;
			25036: outdata = 32'd40500;
			25037: outdata = 32'd40499;
			25038: outdata = 32'd40498;
			25039: outdata = 32'd40497;
			25040: outdata = 32'd40496;
			25041: outdata = 32'd40495;
			25042: outdata = 32'd40494;
			25043: outdata = 32'd40493;
			25044: outdata = 32'd40492;
			25045: outdata = 32'd40491;
			25046: outdata = 32'd40490;
			25047: outdata = 32'd40489;
			25048: outdata = 32'd40488;
			25049: outdata = 32'd40487;
			25050: outdata = 32'd40486;
			25051: outdata = 32'd40485;
			25052: outdata = 32'd40484;
			25053: outdata = 32'd40483;
			25054: outdata = 32'd40482;
			25055: outdata = 32'd40481;
			25056: outdata = 32'd40480;
			25057: outdata = 32'd40479;
			25058: outdata = 32'd40478;
			25059: outdata = 32'd40477;
			25060: outdata = 32'd40476;
			25061: outdata = 32'd40475;
			25062: outdata = 32'd40474;
			25063: outdata = 32'd40473;
			25064: outdata = 32'd40472;
			25065: outdata = 32'd40471;
			25066: outdata = 32'd40470;
			25067: outdata = 32'd40469;
			25068: outdata = 32'd40468;
			25069: outdata = 32'd40467;
			25070: outdata = 32'd40466;
			25071: outdata = 32'd40465;
			25072: outdata = 32'd40464;
			25073: outdata = 32'd40463;
			25074: outdata = 32'd40462;
			25075: outdata = 32'd40461;
			25076: outdata = 32'd40460;
			25077: outdata = 32'd40459;
			25078: outdata = 32'd40458;
			25079: outdata = 32'd40457;
			25080: outdata = 32'd40456;
			25081: outdata = 32'd40455;
			25082: outdata = 32'd40454;
			25083: outdata = 32'd40453;
			25084: outdata = 32'd40452;
			25085: outdata = 32'd40451;
			25086: outdata = 32'd40450;
			25087: outdata = 32'd40449;
			25088: outdata = 32'd40448;
			25089: outdata = 32'd40447;
			25090: outdata = 32'd40446;
			25091: outdata = 32'd40445;
			25092: outdata = 32'd40444;
			25093: outdata = 32'd40443;
			25094: outdata = 32'd40442;
			25095: outdata = 32'd40441;
			25096: outdata = 32'd40440;
			25097: outdata = 32'd40439;
			25098: outdata = 32'd40438;
			25099: outdata = 32'd40437;
			25100: outdata = 32'd40436;
			25101: outdata = 32'd40435;
			25102: outdata = 32'd40434;
			25103: outdata = 32'd40433;
			25104: outdata = 32'd40432;
			25105: outdata = 32'd40431;
			25106: outdata = 32'd40430;
			25107: outdata = 32'd40429;
			25108: outdata = 32'd40428;
			25109: outdata = 32'd40427;
			25110: outdata = 32'd40426;
			25111: outdata = 32'd40425;
			25112: outdata = 32'd40424;
			25113: outdata = 32'd40423;
			25114: outdata = 32'd40422;
			25115: outdata = 32'd40421;
			25116: outdata = 32'd40420;
			25117: outdata = 32'd40419;
			25118: outdata = 32'd40418;
			25119: outdata = 32'd40417;
			25120: outdata = 32'd40416;
			25121: outdata = 32'd40415;
			25122: outdata = 32'd40414;
			25123: outdata = 32'd40413;
			25124: outdata = 32'd40412;
			25125: outdata = 32'd40411;
			25126: outdata = 32'd40410;
			25127: outdata = 32'd40409;
			25128: outdata = 32'd40408;
			25129: outdata = 32'd40407;
			25130: outdata = 32'd40406;
			25131: outdata = 32'd40405;
			25132: outdata = 32'd40404;
			25133: outdata = 32'd40403;
			25134: outdata = 32'd40402;
			25135: outdata = 32'd40401;
			25136: outdata = 32'd40400;
			25137: outdata = 32'd40399;
			25138: outdata = 32'd40398;
			25139: outdata = 32'd40397;
			25140: outdata = 32'd40396;
			25141: outdata = 32'd40395;
			25142: outdata = 32'd40394;
			25143: outdata = 32'd40393;
			25144: outdata = 32'd40392;
			25145: outdata = 32'd40391;
			25146: outdata = 32'd40390;
			25147: outdata = 32'd40389;
			25148: outdata = 32'd40388;
			25149: outdata = 32'd40387;
			25150: outdata = 32'd40386;
			25151: outdata = 32'd40385;
			25152: outdata = 32'd40384;
			25153: outdata = 32'd40383;
			25154: outdata = 32'd40382;
			25155: outdata = 32'd40381;
			25156: outdata = 32'd40380;
			25157: outdata = 32'd40379;
			25158: outdata = 32'd40378;
			25159: outdata = 32'd40377;
			25160: outdata = 32'd40376;
			25161: outdata = 32'd40375;
			25162: outdata = 32'd40374;
			25163: outdata = 32'd40373;
			25164: outdata = 32'd40372;
			25165: outdata = 32'd40371;
			25166: outdata = 32'd40370;
			25167: outdata = 32'd40369;
			25168: outdata = 32'd40368;
			25169: outdata = 32'd40367;
			25170: outdata = 32'd40366;
			25171: outdata = 32'd40365;
			25172: outdata = 32'd40364;
			25173: outdata = 32'd40363;
			25174: outdata = 32'd40362;
			25175: outdata = 32'd40361;
			25176: outdata = 32'd40360;
			25177: outdata = 32'd40359;
			25178: outdata = 32'd40358;
			25179: outdata = 32'd40357;
			25180: outdata = 32'd40356;
			25181: outdata = 32'd40355;
			25182: outdata = 32'd40354;
			25183: outdata = 32'd40353;
			25184: outdata = 32'd40352;
			25185: outdata = 32'd40351;
			25186: outdata = 32'd40350;
			25187: outdata = 32'd40349;
			25188: outdata = 32'd40348;
			25189: outdata = 32'd40347;
			25190: outdata = 32'd40346;
			25191: outdata = 32'd40345;
			25192: outdata = 32'd40344;
			25193: outdata = 32'd40343;
			25194: outdata = 32'd40342;
			25195: outdata = 32'd40341;
			25196: outdata = 32'd40340;
			25197: outdata = 32'd40339;
			25198: outdata = 32'd40338;
			25199: outdata = 32'd40337;
			25200: outdata = 32'd40336;
			25201: outdata = 32'd40335;
			25202: outdata = 32'd40334;
			25203: outdata = 32'd40333;
			25204: outdata = 32'd40332;
			25205: outdata = 32'd40331;
			25206: outdata = 32'd40330;
			25207: outdata = 32'd40329;
			25208: outdata = 32'd40328;
			25209: outdata = 32'd40327;
			25210: outdata = 32'd40326;
			25211: outdata = 32'd40325;
			25212: outdata = 32'd40324;
			25213: outdata = 32'd40323;
			25214: outdata = 32'd40322;
			25215: outdata = 32'd40321;
			25216: outdata = 32'd40320;
			25217: outdata = 32'd40319;
			25218: outdata = 32'd40318;
			25219: outdata = 32'd40317;
			25220: outdata = 32'd40316;
			25221: outdata = 32'd40315;
			25222: outdata = 32'd40314;
			25223: outdata = 32'd40313;
			25224: outdata = 32'd40312;
			25225: outdata = 32'd40311;
			25226: outdata = 32'd40310;
			25227: outdata = 32'd40309;
			25228: outdata = 32'd40308;
			25229: outdata = 32'd40307;
			25230: outdata = 32'd40306;
			25231: outdata = 32'd40305;
			25232: outdata = 32'd40304;
			25233: outdata = 32'd40303;
			25234: outdata = 32'd40302;
			25235: outdata = 32'd40301;
			25236: outdata = 32'd40300;
			25237: outdata = 32'd40299;
			25238: outdata = 32'd40298;
			25239: outdata = 32'd40297;
			25240: outdata = 32'd40296;
			25241: outdata = 32'd40295;
			25242: outdata = 32'd40294;
			25243: outdata = 32'd40293;
			25244: outdata = 32'd40292;
			25245: outdata = 32'd40291;
			25246: outdata = 32'd40290;
			25247: outdata = 32'd40289;
			25248: outdata = 32'd40288;
			25249: outdata = 32'd40287;
			25250: outdata = 32'd40286;
			25251: outdata = 32'd40285;
			25252: outdata = 32'd40284;
			25253: outdata = 32'd40283;
			25254: outdata = 32'd40282;
			25255: outdata = 32'd40281;
			25256: outdata = 32'd40280;
			25257: outdata = 32'd40279;
			25258: outdata = 32'd40278;
			25259: outdata = 32'd40277;
			25260: outdata = 32'd40276;
			25261: outdata = 32'd40275;
			25262: outdata = 32'd40274;
			25263: outdata = 32'd40273;
			25264: outdata = 32'd40272;
			25265: outdata = 32'd40271;
			25266: outdata = 32'd40270;
			25267: outdata = 32'd40269;
			25268: outdata = 32'd40268;
			25269: outdata = 32'd40267;
			25270: outdata = 32'd40266;
			25271: outdata = 32'd40265;
			25272: outdata = 32'd40264;
			25273: outdata = 32'd40263;
			25274: outdata = 32'd40262;
			25275: outdata = 32'd40261;
			25276: outdata = 32'd40260;
			25277: outdata = 32'd40259;
			25278: outdata = 32'd40258;
			25279: outdata = 32'd40257;
			25280: outdata = 32'd40256;
			25281: outdata = 32'd40255;
			25282: outdata = 32'd40254;
			25283: outdata = 32'd40253;
			25284: outdata = 32'd40252;
			25285: outdata = 32'd40251;
			25286: outdata = 32'd40250;
			25287: outdata = 32'd40249;
			25288: outdata = 32'd40248;
			25289: outdata = 32'd40247;
			25290: outdata = 32'd40246;
			25291: outdata = 32'd40245;
			25292: outdata = 32'd40244;
			25293: outdata = 32'd40243;
			25294: outdata = 32'd40242;
			25295: outdata = 32'd40241;
			25296: outdata = 32'd40240;
			25297: outdata = 32'd40239;
			25298: outdata = 32'd40238;
			25299: outdata = 32'd40237;
			25300: outdata = 32'd40236;
			25301: outdata = 32'd40235;
			25302: outdata = 32'd40234;
			25303: outdata = 32'd40233;
			25304: outdata = 32'd40232;
			25305: outdata = 32'd40231;
			25306: outdata = 32'd40230;
			25307: outdata = 32'd40229;
			25308: outdata = 32'd40228;
			25309: outdata = 32'd40227;
			25310: outdata = 32'd40226;
			25311: outdata = 32'd40225;
			25312: outdata = 32'd40224;
			25313: outdata = 32'd40223;
			25314: outdata = 32'd40222;
			25315: outdata = 32'd40221;
			25316: outdata = 32'd40220;
			25317: outdata = 32'd40219;
			25318: outdata = 32'd40218;
			25319: outdata = 32'd40217;
			25320: outdata = 32'd40216;
			25321: outdata = 32'd40215;
			25322: outdata = 32'd40214;
			25323: outdata = 32'd40213;
			25324: outdata = 32'd40212;
			25325: outdata = 32'd40211;
			25326: outdata = 32'd40210;
			25327: outdata = 32'd40209;
			25328: outdata = 32'd40208;
			25329: outdata = 32'd40207;
			25330: outdata = 32'd40206;
			25331: outdata = 32'd40205;
			25332: outdata = 32'd40204;
			25333: outdata = 32'd40203;
			25334: outdata = 32'd40202;
			25335: outdata = 32'd40201;
			25336: outdata = 32'd40200;
			25337: outdata = 32'd40199;
			25338: outdata = 32'd40198;
			25339: outdata = 32'd40197;
			25340: outdata = 32'd40196;
			25341: outdata = 32'd40195;
			25342: outdata = 32'd40194;
			25343: outdata = 32'd40193;
			25344: outdata = 32'd40192;
			25345: outdata = 32'd40191;
			25346: outdata = 32'd40190;
			25347: outdata = 32'd40189;
			25348: outdata = 32'd40188;
			25349: outdata = 32'd40187;
			25350: outdata = 32'd40186;
			25351: outdata = 32'd40185;
			25352: outdata = 32'd40184;
			25353: outdata = 32'd40183;
			25354: outdata = 32'd40182;
			25355: outdata = 32'd40181;
			25356: outdata = 32'd40180;
			25357: outdata = 32'd40179;
			25358: outdata = 32'd40178;
			25359: outdata = 32'd40177;
			25360: outdata = 32'd40176;
			25361: outdata = 32'd40175;
			25362: outdata = 32'd40174;
			25363: outdata = 32'd40173;
			25364: outdata = 32'd40172;
			25365: outdata = 32'd40171;
			25366: outdata = 32'd40170;
			25367: outdata = 32'd40169;
			25368: outdata = 32'd40168;
			25369: outdata = 32'd40167;
			25370: outdata = 32'd40166;
			25371: outdata = 32'd40165;
			25372: outdata = 32'd40164;
			25373: outdata = 32'd40163;
			25374: outdata = 32'd40162;
			25375: outdata = 32'd40161;
			25376: outdata = 32'd40160;
			25377: outdata = 32'd40159;
			25378: outdata = 32'd40158;
			25379: outdata = 32'd40157;
			25380: outdata = 32'd40156;
			25381: outdata = 32'd40155;
			25382: outdata = 32'd40154;
			25383: outdata = 32'd40153;
			25384: outdata = 32'd40152;
			25385: outdata = 32'd40151;
			25386: outdata = 32'd40150;
			25387: outdata = 32'd40149;
			25388: outdata = 32'd40148;
			25389: outdata = 32'd40147;
			25390: outdata = 32'd40146;
			25391: outdata = 32'd40145;
			25392: outdata = 32'd40144;
			25393: outdata = 32'd40143;
			25394: outdata = 32'd40142;
			25395: outdata = 32'd40141;
			25396: outdata = 32'd40140;
			25397: outdata = 32'd40139;
			25398: outdata = 32'd40138;
			25399: outdata = 32'd40137;
			25400: outdata = 32'd40136;
			25401: outdata = 32'd40135;
			25402: outdata = 32'd40134;
			25403: outdata = 32'd40133;
			25404: outdata = 32'd40132;
			25405: outdata = 32'd40131;
			25406: outdata = 32'd40130;
			25407: outdata = 32'd40129;
			25408: outdata = 32'd40128;
			25409: outdata = 32'd40127;
			25410: outdata = 32'd40126;
			25411: outdata = 32'd40125;
			25412: outdata = 32'd40124;
			25413: outdata = 32'd40123;
			25414: outdata = 32'd40122;
			25415: outdata = 32'd40121;
			25416: outdata = 32'd40120;
			25417: outdata = 32'd40119;
			25418: outdata = 32'd40118;
			25419: outdata = 32'd40117;
			25420: outdata = 32'd40116;
			25421: outdata = 32'd40115;
			25422: outdata = 32'd40114;
			25423: outdata = 32'd40113;
			25424: outdata = 32'd40112;
			25425: outdata = 32'd40111;
			25426: outdata = 32'd40110;
			25427: outdata = 32'd40109;
			25428: outdata = 32'd40108;
			25429: outdata = 32'd40107;
			25430: outdata = 32'd40106;
			25431: outdata = 32'd40105;
			25432: outdata = 32'd40104;
			25433: outdata = 32'd40103;
			25434: outdata = 32'd40102;
			25435: outdata = 32'd40101;
			25436: outdata = 32'd40100;
			25437: outdata = 32'd40099;
			25438: outdata = 32'd40098;
			25439: outdata = 32'd40097;
			25440: outdata = 32'd40096;
			25441: outdata = 32'd40095;
			25442: outdata = 32'd40094;
			25443: outdata = 32'd40093;
			25444: outdata = 32'd40092;
			25445: outdata = 32'd40091;
			25446: outdata = 32'd40090;
			25447: outdata = 32'd40089;
			25448: outdata = 32'd40088;
			25449: outdata = 32'd40087;
			25450: outdata = 32'd40086;
			25451: outdata = 32'd40085;
			25452: outdata = 32'd40084;
			25453: outdata = 32'd40083;
			25454: outdata = 32'd40082;
			25455: outdata = 32'd40081;
			25456: outdata = 32'd40080;
			25457: outdata = 32'd40079;
			25458: outdata = 32'd40078;
			25459: outdata = 32'd40077;
			25460: outdata = 32'd40076;
			25461: outdata = 32'd40075;
			25462: outdata = 32'd40074;
			25463: outdata = 32'd40073;
			25464: outdata = 32'd40072;
			25465: outdata = 32'd40071;
			25466: outdata = 32'd40070;
			25467: outdata = 32'd40069;
			25468: outdata = 32'd40068;
			25469: outdata = 32'd40067;
			25470: outdata = 32'd40066;
			25471: outdata = 32'd40065;
			25472: outdata = 32'd40064;
			25473: outdata = 32'd40063;
			25474: outdata = 32'd40062;
			25475: outdata = 32'd40061;
			25476: outdata = 32'd40060;
			25477: outdata = 32'd40059;
			25478: outdata = 32'd40058;
			25479: outdata = 32'd40057;
			25480: outdata = 32'd40056;
			25481: outdata = 32'd40055;
			25482: outdata = 32'd40054;
			25483: outdata = 32'd40053;
			25484: outdata = 32'd40052;
			25485: outdata = 32'd40051;
			25486: outdata = 32'd40050;
			25487: outdata = 32'd40049;
			25488: outdata = 32'd40048;
			25489: outdata = 32'd40047;
			25490: outdata = 32'd40046;
			25491: outdata = 32'd40045;
			25492: outdata = 32'd40044;
			25493: outdata = 32'd40043;
			25494: outdata = 32'd40042;
			25495: outdata = 32'd40041;
			25496: outdata = 32'd40040;
			25497: outdata = 32'd40039;
			25498: outdata = 32'd40038;
			25499: outdata = 32'd40037;
			25500: outdata = 32'd40036;
			25501: outdata = 32'd40035;
			25502: outdata = 32'd40034;
			25503: outdata = 32'd40033;
			25504: outdata = 32'd40032;
			25505: outdata = 32'd40031;
			25506: outdata = 32'd40030;
			25507: outdata = 32'd40029;
			25508: outdata = 32'd40028;
			25509: outdata = 32'd40027;
			25510: outdata = 32'd40026;
			25511: outdata = 32'd40025;
			25512: outdata = 32'd40024;
			25513: outdata = 32'd40023;
			25514: outdata = 32'd40022;
			25515: outdata = 32'd40021;
			25516: outdata = 32'd40020;
			25517: outdata = 32'd40019;
			25518: outdata = 32'd40018;
			25519: outdata = 32'd40017;
			25520: outdata = 32'd40016;
			25521: outdata = 32'd40015;
			25522: outdata = 32'd40014;
			25523: outdata = 32'd40013;
			25524: outdata = 32'd40012;
			25525: outdata = 32'd40011;
			25526: outdata = 32'd40010;
			25527: outdata = 32'd40009;
			25528: outdata = 32'd40008;
			25529: outdata = 32'd40007;
			25530: outdata = 32'd40006;
			25531: outdata = 32'd40005;
			25532: outdata = 32'd40004;
			25533: outdata = 32'd40003;
			25534: outdata = 32'd40002;
			25535: outdata = 32'd40001;
			25536: outdata = 32'd40000;
			25537: outdata = 32'd39999;
			25538: outdata = 32'd39998;
			25539: outdata = 32'd39997;
			25540: outdata = 32'd39996;
			25541: outdata = 32'd39995;
			25542: outdata = 32'd39994;
			25543: outdata = 32'd39993;
			25544: outdata = 32'd39992;
			25545: outdata = 32'd39991;
			25546: outdata = 32'd39990;
			25547: outdata = 32'd39989;
			25548: outdata = 32'd39988;
			25549: outdata = 32'd39987;
			25550: outdata = 32'd39986;
			25551: outdata = 32'd39985;
			25552: outdata = 32'd39984;
			25553: outdata = 32'd39983;
			25554: outdata = 32'd39982;
			25555: outdata = 32'd39981;
			25556: outdata = 32'd39980;
			25557: outdata = 32'd39979;
			25558: outdata = 32'd39978;
			25559: outdata = 32'd39977;
			25560: outdata = 32'd39976;
			25561: outdata = 32'd39975;
			25562: outdata = 32'd39974;
			25563: outdata = 32'd39973;
			25564: outdata = 32'd39972;
			25565: outdata = 32'd39971;
			25566: outdata = 32'd39970;
			25567: outdata = 32'd39969;
			25568: outdata = 32'd39968;
			25569: outdata = 32'd39967;
			25570: outdata = 32'd39966;
			25571: outdata = 32'd39965;
			25572: outdata = 32'd39964;
			25573: outdata = 32'd39963;
			25574: outdata = 32'd39962;
			25575: outdata = 32'd39961;
			25576: outdata = 32'd39960;
			25577: outdata = 32'd39959;
			25578: outdata = 32'd39958;
			25579: outdata = 32'd39957;
			25580: outdata = 32'd39956;
			25581: outdata = 32'd39955;
			25582: outdata = 32'd39954;
			25583: outdata = 32'd39953;
			25584: outdata = 32'd39952;
			25585: outdata = 32'd39951;
			25586: outdata = 32'd39950;
			25587: outdata = 32'd39949;
			25588: outdata = 32'd39948;
			25589: outdata = 32'd39947;
			25590: outdata = 32'd39946;
			25591: outdata = 32'd39945;
			25592: outdata = 32'd39944;
			25593: outdata = 32'd39943;
			25594: outdata = 32'd39942;
			25595: outdata = 32'd39941;
			25596: outdata = 32'd39940;
			25597: outdata = 32'd39939;
			25598: outdata = 32'd39938;
			25599: outdata = 32'd39937;
			25600: outdata = 32'd39936;
			25601: outdata = 32'd39935;
			25602: outdata = 32'd39934;
			25603: outdata = 32'd39933;
			25604: outdata = 32'd39932;
			25605: outdata = 32'd39931;
			25606: outdata = 32'd39930;
			25607: outdata = 32'd39929;
			25608: outdata = 32'd39928;
			25609: outdata = 32'd39927;
			25610: outdata = 32'd39926;
			25611: outdata = 32'd39925;
			25612: outdata = 32'd39924;
			25613: outdata = 32'd39923;
			25614: outdata = 32'd39922;
			25615: outdata = 32'd39921;
			25616: outdata = 32'd39920;
			25617: outdata = 32'd39919;
			25618: outdata = 32'd39918;
			25619: outdata = 32'd39917;
			25620: outdata = 32'd39916;
			25621: outdata = 32'd39915;
			25622: outdata = 32'd39914;
			25623: outdata = 32'd39913;
			25624: outdata = 32'd39912;
			25625: outdata = 32'd39911;
			25626: outdata = 32'd39910;
			25627: outdata = 32'd39909;
			25628: outdata = 32'd39908;
			25629: outdata = 32'd39907;
			25630: outdata = 32'd39906;
			25631: outdata = 32'd39905;
			25632: outdata = 32'd39904;
			25633: outdata = 32'd39903;
			25634: outdata = 32'd39902;
			25635: outdata = 32'd39901;
			25636: outdata = 32'd39900;
			25637: outdata = 32'd39899;
			25638: outdata = 32'd39898;
			25639: outdata = 32'd39897;
			25640: outdata = 32'd39896;
			25641: outdata = 32'd39895;
			25642: outdata = 32'd39894;
			25643: outdata = 32'd39893;
			25644: outdata = 32'd39892;
			25645: outdata = 32'd39891;
			25646: outdata = 32'd39890;
			25647: outdata = 32'd39889;
			25648: outdata = 32'd39888;
			25649: outdata = 32'd39887;
			25650: outdata = 32'd39886;
			25651: outdata = 32'd39885;
			25652: outdata = 32'd39884;
			25653: outdata = 32'd39883;
			25654: outdata = 32'd39882;
			25655: outdata = 32'd39881;
			25656: outdata = 32'd39880;
			25657: outdata = 32'd39879;
			25658: outdata = 32'd39878;
			25659: outdata = 32'd39877;
			25660: outdata = 32'd39876;
			25661: outdata = 32'd39875;
			25662: outdata = 32'd39874;
			25663: outdata = 32'd39873;
			25664: outdata = 32'd39872;
			25665: outdata = 32'd39871;
			25666: outdata = 32'd39870;
			25667: outdata = 32'd39869;
			25668: outdata = 32'd39868;
			25669: outdata = 32'd39867;
			25670: outdata = 32'd39866;
			25671: outdata = 32'd39865;
			25672: outdata = 32'd39864;
			25673: outdata = 32'd39863;
			25674: outdata = 32'd39862;
			25675: outdata = 32'd39861;
			25676: outdata = 32'd39860;
			25677: outdata = 32'd39859;
			25678: outdata = 32'd39858;
			25679: outdata = 32'd39857;
			25680: outdata = 32'd39856;
			25681: outdata = 32'd39855;
			25682: outdata = 32'd39854;
			25683: outdata = 32'd39853;
			25684: outdata = 32'd39852;
			25685: outdata = 32'd39851;
			25686: outdata = 32'd39850;
			25687: outdata = 32'd39849;
			25688: outdata = 32'd39848;
			25689: outdata = 32'd39847;
			25690: outdata = 32'd39846;
			25691: outdata = 32'd39845;
			25692: outdata = 32'd39844;
			25693: outdata = 32'd39843;
			25694: outdata = 32'd39842;
			25695: outdata = 32'd39841;
			25696: outdata = 32'd39840;
			25697: outdata = 32'd39839;
			25698: outdata = 32'd39838;
			25699: outdata = 32'd39837;
			25700: outdata = 32'd39836;
			25701: outdata = 32'd39835;
			25702: outdata = 32'd39834;
			25703: outdata = 32'd39833;
			25704: outdata = 32'd39832;
			25705: outdata = 32'd39831;
			25706: outdata = 32'd39830;
			25707: outdata = 32'd39829;
			25708: outdata = 32'd39828;
			25709: outdata = 32'd39827;
			25710: outdata = 32'd39826;
			25711: outdata = 32'd39825;
			25712: outdata = 32'd39824;
			25713: outdata = 32'd39823;
			25714: outdata = 32'd39822;
			25715: outdata = 32'd39821;
			25716: outdata = 32'd39820;
			25717: outdata = 32'd39819;
			25718: outdata = 32'd39818;
			25719: outdata = 32'd39817;
			25720: outdata = 32'd39816;
			25721: outdata = 32'd39815;
			25722: outdata = 32'd39814;
			25723: outdata = 32'd39813;
			25724: outdata = 32'd39812;
			25725: outdata = 32'd39811;
			25726: outdata = 32'd39810;
			25727: outdata = 32'd39809;
			25728: outdata = 32'd39808;
			25729: outdata = 32'd39807;
			25730: outdata = 32'd39806;
			25731: outdata = 32'd39805;
			25732: outdata = 32'd39804;
			25733: outdata = 32'd39803;
			25734: outdata = 32'd39802;
			25735: outdata = 32'd39801;
			25736: outdata = 32'd39800;
			25737: outdata = 32'd39799;
			25738: outdata = 32'd39798;
			25739: outdata = 32'd39797;
			25740: outdata = 32'd39796;
			25741: outdata = 32'd39795;
			25742: outdata = 32'd39794;
			25743: outdata = 32'd39793;
			25744: outdata = 32'd39792;
			25745: outdata = 32'd39791;
			25746: outdata = 32'd39790;
			25747: outdata = 32'd39789;
			25748: outdata = 32'd39788;
			25749: outdata = 32'd39787;
			25750: outdata = 32'd39786;
			25751: outdata = 32'd39785;
			25752: outdata = 32'd39784;
			25753: outdata = 32'd39783;
			25754: outdata = 32'd39782;
			25755: outdata = 32'd39781;
			25756: outdata = 32'd39780;
			25757: outdata = 32'd39779;
			25758: outdata = 32'd39778;
			25759: outdata = 32'd39777;
			25760: outdata = 32'd39776;
			25761: outdata = 32'd39775;
			25762: outdata = 32'd39774;
			25763: outdata = 32'd39773;
			25764: outdata = 32'd39772;
			25765: outdata = 32'd39771;
			25766: outdata = 32'd39770;
			25767: outdata = 32'd39769;
			25768: outdata = 32'd39768;
			25769: outdata = 32'd39767;
			25770: outdata = 32'd39766;
			25771: outdata = 32'd39765;
			25772: outdata = 32'd39764;
			25773: outdata = 32'd39763;
			25774: outdata = 32'd39762;
			25775: outdata = 32'd39761;
			25776: outdata = 32'd39760;
			25777: outdata = 32'd39759;
			25778: outdata = 32'd39758;
			25779: outdata = 32'd39757;
			25780: outdata = 32'd39756;
			25781: outdata = 32'd39755;
			25782: outdata = 32'd39754;
			25783: outdata = 32'd39753;
			25784: outdata = 32'd39752;
			25785: outdata = 32'd39751;
			25786: outdata = 32'd39750;
			25787: outdata = 32'd39749;
			25788: outdata = 32'd39748;
			25789: outdata = 32'd39747;
			25790: outdata = 32'd39746;
			25791: outdata = 32'd39745;
			25792: outdata = 32'd39744;
			25793: outdata = 32'd39743;
			25794: outdata = 32'd39742;
			25795: outdata = 32'd39741;
			25796: outdata = 32'd39740;
			25797: outdata = 32'd39739;
			25798: outdata = 32'd39738;
			25799: outdata = 32'd39737;
			25800: outdata = 32'd39736;
			25801: outdata = 32'd39735;
			25802: outdata = 32'd39734;
			25803: outdata = 32'd39733;
			25804: outdata = 32'd39732;
			25805: outdata = 32'd39731;
			25806: outdata = 32'd39730;
			25807: outdata = 32'd39729;
			25808: outdata = 32'd39728;
			25809: outdata = 32'd39727;
			25810: outdata = 32'd39726;
			25811: outdata = 32'd39725;
			25812: outdata = 32'd39724;
			25813: outdata = 32'd39723;
			25814: outdata = 32'd39722;
			25815: outdata = 32'd39721;
			25816: outdata = 32'd39720;
			25817: outdata = 32'd39719;
			25818: outdata = 32'd39718;
			25819: outdata = 32'd39717;
			25820: outdata = 32'd39716;
			25821: outdata = 32'd39715;
			25822: outdata = 32'd39714;
			25823: outdata = 32'd39713;
			25824: outdata = 32'd39712;
			25825: outdata = 32'd39711;
			25826: outdata = 32'd39710;
			25827: outdata = 32'd39709;
			25828: outdata = 32'd39708;
			25829: outdata = 32'd39707;
			25830: outdata = 32'd39706;
			25831: outdata = 32'd39705;
			25832: outdata = 32'd39704;
			25833: outdata = 32'd39703;
			25834: outdata = 32'd39702;
			25835: outdata = 32'd39701;
			25836: outdata = 32'd39700;
			25837: outdata = 32'd39699;
			25838: outdata = 32'd39698;
			25839: outdata = 32'd39697;
			25840: outdata = 32'd39696;
			25841: outdata = 32'd39695;
			25842: outdata = 32'd39694;
			25843: outdata = 32'd39693;
			25844: outdata = 32'd39692;
			25845: outdata = 32'd39691;
			25846: outdata = 32'd39690;
			25847: outdata = 32'd39689;
			25848: outdata = 32'd39688;
			25849: outdata = 32'd39687;
			25850: outdata = 32'd39686;
			25851: outdata = 32'd39685;
			25852: outdata = 32'd39684;
			25853: outdata = 32'd39683;
			25854: outdata = 32'd39682;
			25855: outdata = 32'd39681;
			25856: outdata = 32'd39680;
			25857: outdata = 32'd39679;
			25858: outdata = 32'd39678;
			25859: outdata = 32'd39677;
			25860: outdata = 32'd39676;
			25861: outdata = 32'd39675;
			25862: outdata = 32'd39674;
			25863: outdata = 32'd39673;
			25864: outdata = 32'd39672;
			25865: outdata = 32'd39671;
			25866: outdata = 32'd39670;
			25867: outdata = 32'd39669;
			25868: outdata = 32'd39668;
			25869: outdata = 32'd39667;
			25870: outdata = 32'd39666;
			25871: outdata = 32'd39665;
			25872: outdata = 32'd39664;
			25873: outdata = 32'd39663;
			25874: outdata = 32'd39662;
			25875: outdata = 32'd39661;
			25876: outdata = 32'd39660;
			25877: outdata = 32'd39659;
			25878: outdata = 32'd39658;
			25879: outdata = 32'd39657;
			25880: outdata = 32'd39656;
			25881: outdata = 32'd39655;
			25882: outdata = 32'd39654;
			25883: outdata = 32'd39653;
			25884: outdata = 32'd39652;
			25885: outdata = 32'd39651;
			25886: outdata = 32'd39650;
			25887: outdata = 32'd39649;
			25888: outdata = 32'd39648;
			25889: outdata = 32'd39647;
			25890: outdata = 32'd39646;
			25891: outdata = 32'd39645;
			25892: outdata = 32'd39644;
			25893: outdata = 32'd39643;
			25894: outdata = 32'd39642;
			25895: outdata = 32'd39641;
			25896: outdata = 32'd39640;
			25897: outdata = 32'd39639;
			25898: outdata = 32'd39638;
			25899: outdata = 32'd39637;
			25900: outdata = 32'd39636;
			25901: outdata = 32'd39635;
			25902: outdata = 32'd39634;
			25903: outdata = 32'd39633;
			25904: outdata = 32'd39632;
			25905: outdata = 32'd39631;
			25906: outdata = 32'd39630;
			25907: outdata = 32'd39629;
			25908: outdata = 32'd39628;
			25909: outdata = 32'd39627;
			25910: outdata = 32'd39626;
			25911: outdata = 32'd39625;
			25912: outdata = 32'd39624;
			25913: outdata = 32'd39623;
			25914: outdata = 32'd39622;
			25915: outdata = 32'd39621;
			25916: outdata = 32'd39620;
			25917: outdata = 32'd39619;
			25918: outdata = 32'd39618;
			25919: outdata = 32'd39617;
			25920: outdata = 32'd39616;
			25921: outdata = 32'd39615;
			25922: outdata = 32'd39614;
			25923: outdata = 32'd39613;
			25924: outdata = 32'd39612;
			25925: outdata = 32'd39611;
			25926: outdata = 32'd39610;
			25927: outdata = 32'd39609;
			25928: outdata = 32'd39608;
			25929: outdata = 32'd39607;
			25930: outdata = 32'd39606;
			25931: outdata = 32'd39605;
			25932: outdata = 32'd39604;
			25933: outdata = 32'd39603;
			25934: outdata = 32'd39602;
			25935: outdata = 32'd39601;
			25936: outdata = 32'd39600;
			25937: outdata = 32'd39599;
			25938: outdata = 32'd39598;
			25939: outdata = 32'd39597;
			25940: outdata = 32'd39596;
			25941: outdata = 32'd39595;
			25942: outdata = 32'd39594;
			25943: outdata = 32'd39593;
			25944: outdata = 32'd39592;
			25945: outdata = 32'd39591;
			25946: outdata = 32'd39590;
			25947: outdata = 32'd39589;
			25948: outdata = 32'd39588;
			25949: outdata = 32'd39587;
			25950: outdata = 32'd39586;
			25951: outdata = 32'd39585;
			25952: outdata = 32'd39584;
			25953: outdata = 32'd39583;
			25954: outdata = 32'd39582;
			25955: outdata = 32'd39581;
			25956: outdata = 32'd39580;
			25957: outdata = 32'd39579;
			25958: outdata = 32'd39578;
			25959: outdata = 32'd39577;
			25960: outdata = 32'd39576;
			25961: outdata = 32'd39575;
			25962: outdata = 32'd39574;
			25963: outdata = 32'd39573;
			25964: outdata = 32'd39572;
			25965: outdata = 32'd39571;
			25966: outdata = 32'd39570;
			25967: outdata = 32'd39569;
			25968: outdata = 32'd39568;
			25969: outdata = 32'd39567;
			25970: outdata = 32'd39566;
			25971: outdata = 32'd39565;
			25972: outdata = 32'd39564;
			25973: outdata = 32'd39563;
			25974: outdata = 32'd39562;
			25975: outdata = 32'd39561;
			25976: outdata = 32'd39560;
			25977: outdata = 32'd39559;
			25978: outdata = 32'd39558;
			25979: outdata = 32'd39557;
			25980: outdata = 32'd39556;
			25981: outdata = 32'd39555;
			25982: outdata = 32'd39554;
			25983: outdata = 32'd39553;
			25984: outdata = 32'd39552;
			25985: outdata = 32'd39551;
			25986: outdata = 32'd39550;
			25987: outdata = 32'd39549;
			25988: outdata = 32'd39548;
			25989: outdata = 32'd39547;
			25990: outdata = 32'd39546;
			25991: outdata = 32'd39545;
			25992: outdata = 32'd39544;
			25993: outdata = 32'd39543;
			25994: outdata = 32'd39542;
			25995: outdata = 32'd39541;
			25996: outdata = 32'd39540;
			25997: outdata = 32'd39539;
			25998: outdata = 32'd39538;
			25999: outdata = 32'd39537;
			26000: outdata = 32'd39536;
			26001: outdata = 32'd39535;
			26002: outdata = 32'd39534;
			26003: outdata = 32'd39533;
			26004: outdata = 32'd39532;
			26005: outdata = 32'd39531;
			26006: outdata = 32'd39530;
			26007: outdata = 32'd39529;
			26008: outdata = 32'd39528;
			26009: outdata = 32'd39527;
			26010: outdata = 32'd39526;
			26011: outdata = 32'd39525;
			26012: outdata = 32'd39524;
			26013: outdata = 32'd39523;
			26014: outdata = 32'd39522;
			26015: outdata = 32'd39521;
			26016: outdata = 32'd39520;
			26017: outdata = 32'd39519;
			26018: outdata = 32'd39518;
			26019: outdata = 32'd39517;
			26020: outdata = 32'd39516;
			26021: outdata = 32'd39515;
			26022: outdata = 32'd39514;
			26023: outdata = 32'd39513;
			26024: outdata = 32'd39512;
			26025: outdata = 32'd39511;
			26026: outdata = 32'd39510;
			26027: outdata = 32'd39509;
			26028: outdata = 32'd39508;
			26029: outdata = 32'd39507;
			26030: outdata = 32'd39506;
			26031: outdata = 32'd39505;
			26032: outdata = 32'd39504;
			26033: outdata = 32'd39503;
			26034: outdata = 32'd39502;
			26035: outdata = 32'd39501;
			26036: outdata = 32'd39500;
			26037: outdata = 32'd39499;
			26038: outdata = 32'd39498;
			26039: outdata = 32'd39497;
			26040: outdata = 32'd39496;
			26041: outdata = 32'd39495;
			26042: outdata = 32'd39494;
			26043: outdata = 32'd39493;
			26044: outdata = 32'd39492;
			26045: outdata = 32'd39491;
			26046: outdata = 32'd39490;
			26047: outdata = 32'd39489;
			26048: outdata = 32'd39488;
			26049: outdata = 32'd39487;
			26050: outdata = 32'd39486;
			26051: outdata = 32'd39485;
			26052: outdata = 32'd39484;
			26053: outdata = 32'd39483;
			26054: outdata = 32'd39482;
			26055: outdata = 32'd39481;
			26056: outdata = 32'd39480;
			26057: outdata = 32'd39479;
			26058: outdata = 32'd39478;
			26059: outdata = 32'd39477;
			26060: outdata = 32'd39476;
			26061: outdata = 32'd39475;
			26062: outdata = 32'd39474;
			26063: outdata = 32'd39473;
			26064: outdata = 32'd39472;
			26065: outdata = 32'd39471;
			26066: outdata = 32'd39470;
			26067: outdata = 32'd39469;
			26068: outdata = 32'd39468;
			26069: outdata = 32'd39467;
			26070: outdata = 32'd39466;
			26071: outdata = 32'd39465;
			26072: outdata = 32'd39464;
			26073: outdata = 32'd39463;
			26074: outdata = 32'd39462;
			26075: outdata = 32'd39461;
			26076: outdata = 32'd39460;
			26077: outdata = 32'd39459;
			26078: outdata = 32'd39458;
			26079: outdata = 32'd39457;
			26080: outdata = 32'd39456;
			26081: outdata = 32'd39455;
			26082: outdata = 32'd39454;
			26083: outdata = 32'd39453;
			26084: outdata = 32'd39452;
			26085: outdata = 32'd39451;
			26086: outdata = 32'd39450;
			26087: outdata = 32'd39449;
			26088: outdata = 32'd39448;
			26089: outdata = 32'd39447;
			26090: outdata = 32'd39446;
			26091: outdata = 32'd39445;
			26092: outdata = 32'd39444;
			26093: outdata = 32'd39443;
			26094: outdata = 32'd39442;
			26095: outdata = 32'd39441;
			26096: outdata = 32'd39440;
			26097: outdata = 32'd39439;
			26098: outdata = 32'd39438;
			26099: outdata = 32'd39437;
			26100: outdata = 32'd39436;
			26101: outdata = 32'd39435;
			26102: outdata = 32'd39434;
			26103: outdata = 32'd39433;
			26104: outdata = 32'd39432;
			26105: outdata = 32'd39431;
			26106: outdata = 32'd39430;
			26107: outdata = 32'd39429;
			26108: outdata = 32'd39428;
			26109: outdata = 32'd39427;
			26110: outdata = 32'd39426;
			26111: outdata = 32'd39425;
			26112: outdata = 32'd39424;
			26113: outdata = 32'd39423;
			26114: outdata = 32'd39422;
			26115: outdata = 32'd39421;
			26116: outdata = 32'd39420;
			26117: outdata = 32'd39419;
			26118: outdata = 32'd39418;
			26119: outdata = 32'd39417;
			26120: outdata = 32'd39416;
			26121: outdata = 32'd39415;
			26122: outdata = 32'd39414;
			26123: outdata = 32'd39413;
			26124: outdata = 32'd39412;
			26125: outdata = 32'd39411;
			26126: outdata = 32'd39410;
			26127: outdata = 32'd39409;
			26128: outdata = 32'd39408;
			26129: outdata = 32'd39407;
			26130: outdata = 32'd39406;
			26131: outdata = 32'd39405;
			26132: outdata = 32'd39404;
			26133: outdata = 32'd39403;
			26134: outdata = 32'd39402;
			26135: outdata = 32'd39401;
			26136: outdata = 32'd39400;
			26137: outdata = 32'd39399;
			26138: outdata = 32'd39398;
			26139: outdata = 32'd39397;
			26140: outdata = 32'd39396;
			26141: outdata = 32'd39395;
			26142: outdata = 32'd39394;
			26143: outdata = 32'd39393;
			26144: outdata = 32'd39392;
			26145: outdata = 32'd39391;
			26146: outdata = 32'd39390;
			26147: outdata = 32'd39389;
			26148: outdata = 32'd39388;
			26149: outdata = 32'd39387;
			26150: outdata = 32'd39386;
			26151: outdata = 32'd39385;
			26152: outdata = 32'd39384;
			26153: outdata = 32'd39383;
			26154: outdata = 32'd39382;
			26155: outdata = 32'd39381;
			26156: outdata = 32'd39380;
			26157: outdata = 32'd39379;
			26158: outdata = 32'd39378;
			26159: outdata = 32'd39377;
			26160: outdata = 32'd39376;
			26161: outdata = 32'd39375;
			26162: outdata = 32'd39374;
			26163: outdata = 32'd39373;
			26164: outdata = 32'd39372;
			26165: outdata = 32'd39371;
			26166: outdata = 32'd39370;
			26167: outdata = 32'd39369;
			26168: outdata = 32'd39368;
			26169: outdata = 32'd39367;
			26170: outdata = 32'd39366;
			26171: outdata = 32'd39365;
			26172: outdata = 32'd39364;
			26173: outdata = 32'd39363;
			26174: outdata = 32'd39362;
			26175: outdata = 32'd39361;
			26176: outdata = 32'd39360;
			26177: outdata = 32'd39359;
			26178: outdata = 32'd39358;
			26179: outdata = 32'd39357;
			26180: outdata = 32'd39356;
			26181: outdata = 32'd39355;
			26182: outdata = 32'd39354;
			26183: outdata = 32'd39353;
			26184: outdata = 32'd39352;
			26185: outdata = 32'd39351;
			26186: outdata = 32'd39350;
			26187: outdata = 32'd39349;
			26188: outdata = 32'd39348;
			26189: outdata = 32'd39347;
			26190: outdata = 32'd39346;
			26191: outdata = 32'd39345;
			26192: outdata = 32'd39344;
			26193: outdata = 32'd39343;
			26194: outdata = 32'd39342;
			26195: outdata = 32'd39341;
			26196: outdata = 32'd39340;
			26197: outdata = 32'd39339;
			26198: outdata = 32'd39338;
			26199: outdata = 32'd39337;
			26200: outdata = 32'd39336;
			26201: outdata = 32'd39335;
			26202: outdata = 32'd39334;
			26203: outdata = 32'd39333;
			26204: outdata = 32'd39332;
			26205: outdata = 32'd39331;
			26206: outdata = 32'd39330;
			26207: outdata = 32'd39329;
			26208: outdata = 32'd39328;
			26209: outdata = 32'd39327;
			26210: outdata = 32'd39326;
			26211: outdata = 32'd39325;
			26212: outdata = 32'd39324;
			26213: outdata = 32'd39323;
			26214: outdata = 32'd39322;
			26215: outdata = 32'd39321;
			26216: outdata = 32'd39320;
			26217: outdata = 32'd39319;
			26218: outdata = 32'd39318;
			26219: outdata = 32'd39317;
			26220: outdata = 32'd39316;
			26221: outdata = 32'd39315;
			26222: outdata = 32'd39314;
			26223: outdata = 32'd39313;
			26224: outdata = 32'd39312;
			26225: outdata = 32'd39311;
			26226: outdata = 32'd39310;
			26227: outdata = 32'd39309;
			26228: outdata = 32'd39308;
			26229: outdata = 32'd39307;
			26230: outdata = 32'd39306;
			26231: outdata = 32'd39305;
			26232: outdata = 32'd39304;
			26233: outdata = 32'd39303;
			26234: outdata = 32'd39302;
			26235: outdata = 32'd39301;
			26236: outdata = 32'd39300;
			26237: outdata = 32'd39299;
			26238: outdata = 32'd39298;
			26239: outdata = 32'd39297;
			26240: outdata = 32'd39296;
			26241: outdata = 32'd39295;
			26242: outdata = 32'd39294;
			26243: outdata = 32'd39293;
			26244: outdata = 32'd39292;
			26245: outdata = 32'd39291;
			26246: outdata = 32'd39290;
			26247: outdata = 32'd39289;
			26248: outdata = 32'd39288;
			26249: outdata = 32'd39287;
			26250: outdata = 32'd39286;
			26251: outdata = 32'd39285;
			26252: outdata = 32'd39284;
			26253: outdata = 32'd39283;
			26254: outdata = 32'd39282;
			26255: outdata = 32'd39281;
			26256: outdata = 32'd39280;
			26257: outdata = 32'd39279;
			26258: outdata = 32'd39278;
			26259: outdata = 32'd39277;
			26260: outdata = 32'd39276;
			26261: outdata = 32'd39275;
			26262: outdata = 32'd39274;
			26263: outdata = 32'd39273;
			26264: outdata = 32'd39272;
			26265: outdata = 32'd39271;
			26266: outdata = 32'd39270;
			26267: outdata = 32'd39269;
			26268: outdata = 32'd39268;
			26269: outdata = 32'd39267;
			26270: outdata = 32'd39266;
			26271: outdata = 32'd39265;
			26272: outdata = 32'd39264;
			26273: outdata = 32'd39263;
			26274: outdata = 32'd39262;
			26275: outdata = 32'd39261;
			26276: outdata = 32'd39260;
			26277: outdata = 32'd39259;
			26278: outdata = 32'd39258;
			26279: outdata = 32'd39257;
			26280: outdata = 32'd39256;
			26281: outdata = 32'd39255;
			26282: outdata = 32'd39254;
			26283: outdata = 32'd39253;
			26284: outdata = 32'd39252;
			26285: outdata = 32'd39251;
			26286: outdata = 32'd39250;
			26287: outdata = 32'd39249;
			26288: outdata = 32'd39248;
			26289: outdata = 32'd39247;
			26290: outdata = 32'd39246;
			26291: outdata = 32'd39245;
			26292: outdata = 32'd39244;
			26293: outdata = 32'd39243;
			26294: outdata = 32'd39242;
			26295: outdata = 32'd39241;
			26296: outdata = 32'd39240;
			26297: outdata = 32'd39239;
			26298: outdata = 32'd39238;
			26299: outdata = 32'd39237;
			26300: outdata = 32'd39236;
			26301: outdata = 32'd39235;
			26302: outdata = 32'd39234;
			26303: outdata = 32'd39233;
			26304: outdata = 32'd39232;
			26305: outdata = 32'd39231;
			26306: outdata = 32'd39230;
			26307: outdata = 32'd39229;
			26308: outdata = 32'd39228;
			26309: outdata = 32'd39227;
			26310: outdata = 32'd39226;
			26311: outdata = 32'd39225;
			26312: outdata = 32'd39224;
			26313: outdata = 32'd39223;
			26314: outdata = 32'd39222;
			26315: outdata = 32'd39221;
			26316: outdata = 32'd39220;
			26317: outdata = 32'd39219;
			26318: outdata = 32'd39218;
			26319: outdata = 32'd39217;
			26320: outdata = 32'd39216;
			26321: outdata = 32'd39215;
			26322: outdata = 32'd39214;
			26323: outdata = 32'd39213;
			26324: outdata = 32'd39212;
			26325: outdata = 32'd39211;
			26326: outdata = 32'd39210;
			26327: outdata = 32'd39209;
			26328: outdata = 32'd39208;
			26329: outdata = 32'd39207;
			26330: outdata = 32'd39206;
			26331: outdata = 32'd39205;
			26332: outdata = 32'd39204;
			26333: outdata = 32'd39203;
			26334: outdata = 32'd39202;
			26335: outdata = 32'd39201;
			26336: outdata = 32'd39200;
			26337: outdata = 32'd39199;
			26338: outdata = 32'd39198;
			26339: outdata = 32'd39197;
			26340: outdata = 32'd39196;
			26341: outdata = 32'd39195;
			26342: outdata = 32'd39194;
			26343: outdata = 32'd39193;
			26344: outdata = 32'd39192;
			26345: outdata = 32'd39191;
			26346: outdata = 32'd39190;
			26347: outdata = 32'd39189;
			26348: outdata = 32'd39188;
			26349: outdata = 32'd39187;
			26350: outdata = 32'd39186;
			26351: outdata = 32'd39185;
			26352: outdata = 32'd39184;
			26353: outdata = 32'd39183;
			26354: outdata = 32'd39182;
			26355: outdata = 32'd39181;
			26356: outdata = 32'd39180;
			26357: outdata = 32'd39179;
			26358: outdata = 32'd39178;
			26359: outdata = 32'd39177;
			26360: outdata = 32'd39176;
			26361: outdata = 32'd39175;
			26362: outdata = 32'd39174;
			26363: outdata = 32'd39173;
			26364: outdata = 32'd39172;
			26365: outdata = 32'd39171;
			26366: outdata = 32'd39170;
			26367: outdata = 32'd39169;
			26368: outdata = 32'd39168;
			26369: outdata = 32'd39167;
			26370: outdata = 32'd39166;
			26371: outdata = 32'd39165;
			26372: outdata = 32'd39164;
			26373: outdata = 32'd39163;
			26374: outdata = 32'd39162;
			26375: outdata = 32'd39161;
			26376: outdata = 32'd39160;
			26377: outdata = 32'd39159;
			26378: outdata = 32'd39158;
			26379: outdata = 32'd39157;
			26380: outdata = 32'd39156;
			26381: outdata = 32'd39155;
			26382: outdata = 32'd39154;
			26383: outdata = 32'd39153;
			26384: outdata = 32'd39152;
			26385: outdata = 32'd39151;
			26386: outdata = 32'd39150;
			26387: outdata = 32'd39149;
			26388: outdata = 32'd39148;
			26389: outdata = 32'd39147;
			26390: outdata = 32'd39146;
			26391: outdata = 32'd39145;
			26392: outdata = 32'd39144;
			26393: outdata = 32'd39143;
			26394: outdata = 32'd39142;
			26395: outdata = 32'd39141;
			26396: outdata = 32'd39140;
			26397: outdata = 32'd39139;
			26398: outdata = 32'd39138;
			26399: outdata = 32'd39137;
			26400: outdata = 32'd39136;
			26401: outdata = 32'd39135;
			26402: outdata = 32'd39134;
			26403: outdata = 32'd39133;
			26404: outdata = 32'd39132;
			26405: outdata = 32'd39131;
			26406: outdata = 32'd39130;
			26407: outdata = 32'd39129;
			26408: outdata = 32'd39128;
			26409: outdata = 32'd39127;
			26410: outdata = 32'd39126;
			26411: outdata = 32'd39125;
			26412: outdata = 32'd39124;
			26413: outdata = 32'd39123;
			26414: outdata = 32'd39122;
			26415: outdata = 32'd39121;
			26416: outdata = 32'd39120;
			26417: outdata = 32'd39119;
			26418: outdata = 32'd39118;
			26419: outdata = 32'd39117;
			26420: outdata = 32'd39116;
			26421: outdata = 32'd39115;
			26422: outdata = 32'd39114;
			26423: outdata = 32'd39113;
			26424: outdata = 32'd39112;
			26425: outdata = 32'd39111;
			26426: outdata = 32'd39110;
			26427: outdata = 32'd39109;
			26428: outdata = 32'd39108;
			26429: outdata = 32'd39107;
			26430: outdata = 32'd39106;
			26431: outdata = 32'd39105;
			26432: outdata = 32'd39104;
			26433: outdata = 32'd39103;
			26434: outdata = 32'd39102;
			26435: outdata = 32'd39101;
			26436: outdata = 32'd39100;
			26437: outdata = 32'd39099;
			26438: outdata = 32'd39098;
			26439: outdata = 32'd39097;
			26440: outdata = 32'd39096;
			26441: outdata = 32'd39095;
			26442: outdata = 32'd39094;
			26443: outdata = 32'd39093;
			26444: outdata = 32'd39092;
			26445: outdata = 32'd39091;
			26446: outdata = 32'd39090;
			26447: outdata = 32'd39089;
			26448: outdata = 32'd39088;
			26449: outdata = 32'd39087;
			26450: outdata = 32'd39086;
			26451: outdata = 32'd39085;
			26452: outdata = 32'd39084;
			26453: outdata = 32'd39083;
			26454: outdata = 32'd39082;
			26455: outdata = 32'd39081;
			26456: outdata = 32'd39080;
			26457: outdata = 32'd39079;
			26458: outdata = 32'd39078;
			26459: outdata = 32'd39077;
			26460: outdata = 32'd39076;
			26461: outdata = 32'd39075;
			26462: outdata = 32'd39074;
			26463: outdata = 32'd39073;
			26464: outdata = 32'd39072;
			26465: outdata = 32'd39071;
			26466: outdata = 32'd39070;
			26467: outdata = 32'd39069;
			26468: outdata = 32'd39068;
			26469: outdata = 32'd39067;
			26470: outdata = 32'd39066;
			26471: outdata = 32'd39065;
			26472: outdata = 32'd39064;
			26473: outdata = 32'd39063;
			26474: outdata = 32'd39062;
			26475: outdata = 32'd39061;
			26476: outdata = 32'd39060;
			26477: outdata = 32'd39059;
			26478: outdata = 32'd39058;
			26479: outdata = 32'd39057;
			26480: outdata = 32'd39056;
			26481: outdata = 32'd39055;
			26482: outdata = 32'd39054;
			26483: outdata = 32'd39053;
			26484: outdata = 32'd39052;
			26485: outdata = 32'd39051;
			26486: outdata = 32'd39050;
			26487: outdata = 32'd39049;
			26488: outdata = 32'd39048;
			26489: outdata = 32'd39047;
			26490: outdata = 32'd39046;
			26491: outdata = 32'd39045;
			26492: outdata = 32'd39044;
			26493: outdata = 32'd39043;
			26494: outdata = 32'd39042;
			26495: outdata = 32'd39041;
			26496: outdata = 32'd39040;
			26497: outdata = 32'd39039;
			26498: outdata = 32'd39038;
			26499: outdata = 32'd39037;
			26500: outdata = 32'd39036;
			26501: outdata = 32'd39035;
			26502: outdata = 32'd39034;
			26503: outdata = 32'd39033;
			26504: outdata = 32'd39032;
			26505: outdata = 32'd39031;
			26506: outdata = 32'd39030;
			26507: outdata = 32'd39029;
			26508: outdata = 32'd39028;
			26509: outdata = 32'd39027;
			26510: outdata = 32'd39026;
			26511: outdata = 32'd39025;
			26512: outdata = 32'd39024;
			26513: outdata = 32'd39023;
			26514: outdata = 32'd39022;
			26515: outdata = 32'd39021;
			26516: outdata = 32'd39020;
			26517: outdata = 32'd39019;
			26518: outdata = 32'd39018;
			26519: outdata = 32'd39017;
			26520: outdata = 32'd39016;
			26521: outdata = 32'd39015;
			26522: outdata = 32'd39014;
			26523: outdata = 32'd39013;
			26524: outdata = 32'd39012;
			26525: outdata = 32'd39011;
			26526: outdata = 32'd39010;
			26527: outdata = 32'd39009;
			26528: outdata = 32'd39008;
			26529: outdata = 32'd39007;
			26530: outdata = 32'd39006;
			26531: outdata = 32'd39005;
			26532: outdata = 32'd39004;
			26533: outdata = 32'd39003;
			26534: outdata = 32'd39002;
			26535: outdata = 32'd39001;
			26536: outdata = 32'd39000;
			26537: outdata = 32'd38999;
			26538: outdata = 32'd38998;
			26539: outdata = 32'd38997;
			26540: outdata = 32'd38996;
			26541: outdata = 32'd38995;
			26542: outdata = 32'd38994;
			26543: outdata = 32'd38993;
			26544: outdata = 32'd38992;
			26545: outdata = 32'd38991;
			26546: outdata = 32'd38990;
			26547: outdata = 32'd38989;
			26548: outdata = 32'd38988;
			26549: outdata = 32'd38987;
			26550: outdata = 32'd38986;
			26551: outdata = 32'd38985;
			26552: outdata = 32'd38984;
			26553: outdata = 32'd38983;
			26554: outdata = 32'd38982;
			26555: outdata = 32'd38981;
			26556: outdata = 32'd38980;
			26557: outdata = 32'd38979;
			26558: outdata = 32'd38978;
			26559: outdata = 32'd38977;
			26560: outdata = 32'd38976;
			26561: outdata = 32'd38975;
			26562: outdata = 32'd38974;
			26563: outdata = 32'd38973;
			26564: outdata = 32'd38972;
			26565: outdata = 32'd38971;
			26566: outdata = 32'd38970;
			26567: outdata = 32'd38969;
			26568: outdata = 32'd38968;
			26569: outdata = 32'd38967;
			26570: outdata = 32'd38966;
			26571: outdata = 32'd38965;
			26572: outdata = 32'd38964;
			26573: outdata = 32'd38963;
			26574: outdata = 32'd38962;
			26575: outdata = 32'd38961;
			26576: outdata = 32'd38960;
			26577: outdata = 32'd38959;
			26578: outdata = 32'd38958;
			26579: outdata = 32'd38957;
			26580: outdata = 32'd38956;
			26581: outdata = 32'd38955;
			26582: outdata = 32'd38954;
			26583: outdata = 32'd38953;
			26584: outdata = 32'd38952;
			26585: outdata = 32'd38951;
			26586: outdata = 32'd38950;
			26587: outdata = 32'd38949;
			26588: outdata = 32'd38948;
			26589: outdata = 32'd38947;
			26590: outdata = 32'd38946;
			26591: outdata = 32'd38945;
			26592: outdata = 32'd38944;
			26593: outdata = 32'd38943;
			26594: outdata = 32'd38942;
			26595: outdata = 32'd38941;
			26596: outdata = 32'd38940;
			26597: outdata = 32'd38939;
			26598: outdata = 32'd38938;
			26599: outdata = 32'd38937;
			26600: outdata = 32'd38936;
			26601: outdata = 32'd38935;
			26602: outdata = 32'd38934;
			26603: outdata = 32'd38933;
			26604: outdata = 32'd38932;
			26605: outdata = 32'd38931;
			26606: outdata = 32'd38930;
			26607: outdata = 32'd38929;
			26608: outdata = 32'd38928;
			26609: outdata = 32'd38927;
			26610: outdata = 32'd38926;
			26611: outdata = 32'd38925;
			26612: outdata = 32'd38924;
			26613: outdata = 32'd38923;
			26614: outdata = 32'd38922;
			26615: outdata = 32'd38921;
			26616: outdata = 32'd38920;
			26617: outdata = 32'd38919;
			26618: outdata = 32'd38918;
			26619: outdata = 32'd38917;
			26620: outdata = 32'd38916;
			26621: outdata = 32'd38915;
			26622: outdata = 32'd38914;
			26623: outdata = 32'd38913;
			26624: outdata = 32'd38912;
			26625: outdata = 32'd38911;
			26626: outdata = 32'd38910;
			26627: outdata = 32'd38909;
			26628: outdata = 32'd38908;
			26629: outdata = 32'd38907;
			26630: outdata = 32'd38906;
			26631: outdata = 32'd38905;
			26632: outdata = 32'd38904;
			26633: outdata = 32'd38903;
			26634: outdata = 32'd38902;
			26635: outdata = 32'd38901;
			26636: outdata = 32'd38900;
			26637: outdata = 32'd38899;
			26638: outdata = 32'd38898;
			26639: outdata = 32'd38897;
			26640: outdata = 32'd38896;
			26641: outdata = 32'd38895;
			26642: outdata = 32'd38894;
			26643: outdata = 32'd38893;
			26644: outdata = 32'd38892;
			26645: outdata = 32'd38891;
			26646: outdata = 32'd38890;
			26647: outdata = 32'd38889;
			26648: outdata = 32'd38888;
			26649: outdata = 32'd38887;
			26650: outdata = 32'd38886;
			26651: outdata = 32'd38885;
			26652: outdata = 32'd38884;
			26653: outdata = 32'd38883;
			26654: outdata = 32'd38882;
			26655: outdata = 32'd38881;
			26656: outdata = 32'd38880;
			26657: outdata = 32'd38879;
			26658: outdata = 32'd38878;
			26659: outdata = 32'd38877;
			26660: outdata = 32'd38876;
			26661: outdata = 32'd38875;
			26662: outdata = 32'd38874;
			26663: outdata = 32'd38873;
			26664: outdata = 32'd38872;
			26665: outdata = 32'd38871;
			26666: outdata = 32'd38870;
			26667: outdata = 32'd38869;
			26668: outdata = 32'd38868;
			26669: outdata = 32'd38867;
			26670: outdata = 32'd38866;
			26671: outdata = 32'd38865;
			26672: outdata = 32'd38864;
			26673: outdata = 32'd38863;
			26674: outdata = 32'd38862;
			26675: outdata = 32'd38861;
			26676: outdata = 32'd38860;
			26677: outdata = 32'd38859;
			26678: outdata = 32'd38858;
			26679: outdata = 32'd38857;
			26680: outdata = 32'd38856;
			26681: outdata = 32'd38855;
			26682: outdata = 32'd38854;
			26683: outdata = 32'd38853;
			26684: outdata = 32'd38852;
			26685: outdata = 32'd38851;
			26686: outdata = 32'd38850;
			26687: outdata = 32'd38849;
			26688: outdata = 32'd38848;
			26689: outdata = 32'd38847;
			26690: outdata = 32'd38846;
			26691: outdata = 32'd38845;
			26692: outdata = 32'd38844;
			26693: outdata = 32'd38843;
			26694: outdata = 32'd38842;
			26695: outdata = 32'd38841;
			26696: outdata = 32'd38840;
			26697: outdata = 32'd38839;
			26698: outdata = 32'd38838;
			26699: outdata = 32'd38837;
			26700: outdata = 32'd38836;
			26701: outdata = 32'd38835;
			26702: outdata = 32'd38834;
			26703: outdata = 32'd38833;
			26704: outdata = 32'd38832;
			26705: outdata = 32'd38831;
			26706: outdata = 32'd38830;
			26707: outdata = 32'd38829;
			26708: outdata = 32'd38828;
			26709: outdata = 32'd38827;
			26710: outdata = 32'd38826;
			26711: outdata = 32'd38825;
			26712: outdata = 32'd38824;
			26713: outdata = 32'd38823;
			26714: outdata = 32'd38822;
			26715: outdata = 32'd38821;
			26716: outdata = 32'd38820;
			26717: outdata = 32'd38819;
			26718: outdata = 32'd38818;
			26719: outdata = 32'd38817;
			26720: outdata = 32'd38816;
			26721: outdata = 32'd38815;
			26722: outdata = 32'd38814;
			26723: outdata = 32'd38813;
			26724: outdata = 32'd38812;
			26725: outdata = 32'd38811;
			26726: outdata = 32'd38810;
			26727: outdata = 32'd38809;
			26728: outdata = 32'd38808;
			26729: outdata = 32'd38807;
			26730: outdata = 32'd38806;
			26731: outdata = 32'd38805;
			26732: outdata = 32'd38804;
			26733: outdata = 32'd38803;
			26734: outdata = 32'd38802;
			26735: outdata = 32'd38801;
			26736: outdata = 32'd38800;
			26737: outdata = 32'd38799;
			26738: outdata = 32'd38798;
			26739: outdata = 32'd38797;
			26740: outdata = 32'd38796;
			26741: outdata = 32'd38795;
			26742: outdata = 32'd38794;
			26743: outdata = 32'd38793;
			26744: outdata = 32'd38792;
			26745: outdata = 32'd38791;
			26746: outdata = 32'd38790;
			26747: outdata = 32'd38789;
			26748: outdata = 32'd38788;
			26749: outdata = 32'd38787;
			26750: outdata = 32'd38786;
			26751: outdata = 32'd38785;
			26752: outdata = 32'd38784;
			26753: outdata = 32'd38783;
			26754: outdata = 32'd38782;
			26755: outdata = 32'd38781;
			26756: outdata = 32'd38780;
			26757: outdata = 32'd38779;
			26758: outdata = 32'd38778;
			26759: outdata = 32'd38777;
			26760: outdata = 32'd38776;
			26761: outdata = 32'd38775;
			26762: outdata = 32'd38774;
			26763: outdata = 32'd38773;
			26764: outdata = 32'd38772;
			26765: outdata = 32'd38771;
			26766: outdata = 32'd38770;
			26767: outdata = 32'd38769;
			26768: outdata = 32'd38768;
			26769: outdata = 32'd38767;
			26770: outdata = 32'd38766;
			26771: outdata = 32'd38765;
			26772: outdata = 32'd38764;
			26773: outdata = 32'd38763;
			26774: outdata = 32'd38762;
			26775: outdata = 32'd38761;
			26776: outdata = 32'd38760;
			26777: outdata = 32'd38759;
			26778: outdata = 32'd38758;
			26779: outdata = 32'd38757;
			26780: outdata = 32'd38756;
			26781: outdata = 32'd38755;
			26782: outdata = 32'd38754;
			26783: outdata = 32'd38753;
			26784: outdata = 32'd38752;
			26785: outdata = 32'd38751;
			26786: outdata = 32'd38750;
			26787: outdata = 32'd38749;
			26788: outdata = 32'd38748;
			26789: outdata = 32'd38747;
			26790: outdata = 32'd38746;
			26791: outdata = 32'd38745;
			26792: outdata = 32'd38744;
			26793: outdata = 32'd38743;
			26794: outdata = 32'd38742;
			26795: outdata = 32'd38741;
			26796: outdata = 32'd38740;
			26797: outdata = 32'd38739;
			26798: outdata = 32'd38738;
			26799: outdata = 32'd38737;
			26800: outdata = 32'd38736;
			26801: outdata = 32'd38735;
			26802: outdata = 32'd38734;
			26803: outdata = 32'd38733;
			26804: outdata = 32'd38732;
			26805: outdata = 32'd38731;
			26806: outdata = 32'd38730;
			26807: outdata = 32'd38729;
			26808: outdata = 32'd38728;
			26809: outdata = 32'd38727;
			26810: outdata = 32'd38726;
			26811: outdata = 32'd38725;
			26812: outdata = 32'd38724;
			26813: outdata = 32'd38723;
			26814: outdata = 32'd38722;
			26815: outdata = 32'd38721;
			26816: outdata = 32'd38720;
			26817: outdata = 32'd38719;
			26818: outdata = 32'd38718;
			26819: outdata = 32'd38717;
			26820: outdata = 32'd38716;
			26821: outdata = 32'd38715;
			26822: outdata = 32'd38714;
			26823: outdata = 32'd38713;
			26824: outdata = 32'd38712;
			26825: outdata = 32'd38711;
			26826: outdata = 32'd38710;
			26827: outdata = 32'd38709;
			26828: outdata = 32'd38708;
			26829: outdata = 32'd38707;
			26830: outdata = 32'd38706;
			26831: outdata = 32'd38705;
			26832: outdata = 32'd38704;
			26833: outdata = 32'd38703;
			26834: outdata = 32'd38702;
			26835: outdata = 32'd38701;
			26836: outdata = 32'd38700;
			26837: outdata = 32'd38699;
			26838: outdata = 32'd38698;
			26839: outdata = 32'd38697;
			26840: outdata = 32'd38696;
			26841: outdata = 32'd38695;
			26842: outdata = 32'd38694;
			26843: outdata = 32'd38693;
			26844: outdata = 32'd38692;
			26845: outdata = 32'd38691;
			26846: outdata = 32'd38690;
			26847: outdata = 32'd38689;
			26848: outdata = 32'd38688;
			26849: outdata = 32'd38687;
			26850: outdata = 32'd38686;
			26851: outdata = 32'd38685;
			26852: outdata = 32'd38684;
			26853: outdata = 32'd38683;
			26854: outdata = 32'd38682;
			26855: outdata = 32'd38681;
			26856: outdata = 32'd38680;
			26857: outdata = 32'd38679;
			26858: outdata = 32'd38678;
			26859: outdata = 32'd38677;
			26860: outdata = 32'd38676;
			26861: outdata = 32'd38675;
			26862: outdata = 32'd38674;
			26863: outdata = 32'd38673;
			26864: outdata = 32'd38672;
			26865: outdata = 32'd38671;
			26866: outdata = 32'd38670;
			26867: outdata = 32'd38669;
			26868: outdata = 32'd38668;
			26869: outdata = 32'd38667;
			26870: outdata = 32'd38666;
			26871: outdata = 32'd38665;
			26872: outdata = 32'd38664;
			26873: outdata = 32'd38663;
			26874: outdata = 32'd38662;
			26875: outdata = 32'd38661;
			26876: outdata = 32'd38660;
			26877: outdata = 32'd38659;
			26878: outdata = 32'd38658;
			26879: outdata = 32'd38657;
			26880: outdata = 32'd38656;
			26881: outdata = 32'd38655;
			26882: outdata = 32'd38654;
			26883: outdata = 32'd38653;
			26884: outdata = 32'd38652;
			26885: outdata = 32'd38651;
			26886: outdata = 32'd38650;
			26887: outdata = 32'd38649;
			26888: outdata = 32'd38648;
			26889: outdata = 32'd38647;
			26890: outdata = 32'd38646;
			26891: outdata = 32'd38645;
			26892: outdata = 32'd38644;
			26893: outdata = 32'd38643;
			26894: outdata = 32'd38642;
			26895: outdata = 32'd38641;
			26896: outdata = 32'd38640;
			26897: outdata = 32'd38639;
			26898: outdata = 32'd38638;
			26899: outdata = 32'd38637;
			26900: outdata = 32'd38636;
			26901: outdata = 32'd38635;
			26902: outdata = 32'd38634;
			26903: outdata = 32'd38633;
			26904: outdata = 32'd38632;
			26905: outdata = 32'd38631;
			26906: outdata = 32'd38630;
			26907: outdata = 32'd38629;
			26908: outdata = 32'd38628;
			26909: outdata = 32'd38627;
			26910: outdata = 32'd38626;
			26911: outdata = 32'd38625;
			26912: outdata = 32'd38624;
			26913: outdata = 32'd38623;
			26914: outdata = 32'd38622;
			26915: outdata = 32'd38621;
			26916: outdata = 32'd38620;
			26917: outdata = 32'd38619;
			26918: outdata = 32'd38618;
			26919: outdata = 32'd38617;
			26920: outdata = 32'd38616;
			26921: outdata = 32'd38615;
			26922: outdata = 32'd38614;
			26923: outdata = 32'd38613;
			26924: outdata = 32'd38612;
			26925: outdata = 32'd38611;
			26926: outdata = 32'd38610;
			26927: outdata = 32'd38609;
			26928: outdata = 32'd38608;
			26929: outdata = 32'd38607;
			26930: outdata = 32'd38606;
			26931: outdata = 32'd38605;
			26932: outdata = 32'd38604;
			26933: outdata = 32'd38603;
			26934: outdata = 32'd38602;
			26935: outdata = 32'd38601;
			26936: outdata = 32'd38600;
			26937: outdata = 32'd38599;
			26938: outdata = 32'd38598;
			26939: outdata = 32'd38597;
			26940: outdata = 32'd38596;
			26941: outdata = 32'd38595;
			26942: outdata = 32'd38594;
			26943: outdata = 32'd38593;
			26944: outdata = 32'd38592;
			26945: outdata = 32'd38591;
			26946: outdata = 32'd38590;
			26947: outdata = 32'd38589;
			26948: outdata = 32'd38588;
			26949: outdata = 32'd38587;
			26950: outdata = 32'd38586;
			26951: outdata = 32'd38585;
			26952: outdata = 32'd38584;
			26953: outdata = 32'd38583;
			26954: outdata = 32'd38582;
			26955: outdata = 32'd38581;
			26956: outdata = 32'd38580;
			26957: outdata = 32'd38579;
			26958: outdata = 32'd38578;
			26959: outdata = 32'd38577;
			26960: outdata = 32'd38576;
			26961: outdata = 32'd38575;
			26962: outdata = 32'd38574;
			26963: outdata = 32'd38573;
			26964: outdata = 32'd38572;
			26965: outdata = 32'd38571;
			26966: outdata = 32'd38570;
			26967: outdata = 32'd38569;
			26968: outdata = 32'd38568;
			26969: outdata = 32'd38567;
			26970: outdata = 32'd38566;
			26971: outdata = 32'd38565;
			26972: outdata = 32'd38564;
			26973: outdata = 32'd38563;
			26974: outdata = 32'd38562;
			26975: outdata = 32'd38561;
			26976: outdata = 32'd38560;
			26977: outdata = 32'd38559;
			26978: outdata = 32'd38558;
			26979: outdata = 32'd38557;
			26980: outdata = 32'd38556;
			26981: outdata = 32'd38555;
			26982: outdata = 32'd38554;
			26983: outdata = 32'd38553;
			26984: outdata = 32'd38552;
			26985: outdata = 32'd38551;
			26986: outdata = 32'd38550;
			26987: outdata = 32'd38549;
			26988: outdata = 32'd38548;
			26989: outdata = 32'd38547;
			26990: outdata = 32'd38546;
			26991: outdata = 32'd38545;
			26992: outdata = 32'd38544;
			26993: outdata = 32'd38543;
			26994: outdata = 32'd38542;
			26995: outdata = 32'd38541;
			26996: outdata = 32'd38540;
			26997: outdata = 32'd38539;
			26998: outdata = 32'd38538;
			26999: outdata = 32'd38537;
			27000: outdata = 32'd38536;
			27001: outdata = 32'd38535;
			27002: outdata = 32'd38534;
			27003: outdata = 32'd38533;
			27004: outdata = 32'd38532;
			27005: outdata = 32'd38531;
			27006: outdata = 32'd38530;
			27007: outdata = 32'd38529;
			27008: outdata = 32'd38528;
			27009: outdata = 32'd38527;
			27010: outdata = 32'd38526;
			27011: outdata = 32'd38525;
			27012: outdata = 32'd38524;
			27013: outdata = 32'd38523;
			27014: outdata = 32'd38522;
			27015: outdata = 32'd38521;
			27016: outdata = 32'd38520;
			27017: outdata = 32'd38519;
			27018: outdata = 32'd38518;
			27019: outdata = 32'd38517;
			27020: outdata = 32'd38516;
			27021: outdata = 32'd38515;
			27022: outdata = 32'd38514;
			27023: outdata = 32'd38513;
			27024: outdata = 32'd38512;
			27025: outdata = 32'd38511;
			27026: outdata = 32'd38510;
			27027: outdata = 32'd38509;
			27028: outdata = 32'd38508;
			27029: outdata = 32'd38507;
			27030: outdata = 32'd38506;
			27031: outdata = 32'd38505;
			27032: outdata = 32'd38504;
			27033: outdata = 32'd38503;
			27034: outdata = 32'd38502;
			27035: outdata = 32'd38501;
			27036: outdata = 32'd38500;
			27037: outdata = 32'd38499;
			27038: outdata = 32'd38498;
			27039: outdata = 32'd38497;
			27040: outdata = 32'd38496;
			27041: outdata = 32'd38495;
			27042: outdata = 32'd38494;
			27043: outdata = 32'd38493;
			27044: outdata = 32'd38492;
			27045: outdata = 32'd38491;
			27046: outdata = 32'd38490;
			27047: outdata = 32'd38489;
			27048: outdata = 32'd38488;
			27049: outdata = 32'd38487;
			27050: outdata = 32'd38486;
			27051: outdata = 32'd38485;
			27052: outdata = 32'd38484;
			27053: outdata = 32'd38483;
			27054: outdata = 32'd38482;
			27055: outdata = 32'd38481;
			27056: outdata = 32'd38480;
			27057: outdata = 32'd38479;
			27058: outdata = 32'd38478;
			27059: outdata = 32'd38477;
			27060: outdata = 32'd38476;
			27061: outdata = 32'd38475;
			27062: outdata = 32'd38474;
			27063: outdata = 32'd38473;
			27064: outdata = 32'd38472;
			27065: outdata = 32'd38471;
			27066: outdata = 32'd38470;
			27067: outdata = 32'd38469;
			27068: outdata = 32'd38468;
			27069: outdata = 32'd38467;
			27070: outdata = 32'd38466;
			27071: outdata = 32'd38465;
			27072: outdata = 32'd38464;
			27073: outdata = 32'd38463;
			27074: outdata = 32'd38462;
			27075: outdata = 32'd38461;
			27076: outdata = 32'd38460;
			27077: outdata = 32'd38459;
			27078: outdata = 32'd38458;
			27079: outdata = 32'd38457;
			27080: outdata = 32'd38456;
			27081: outdata = 32'd38455;
			27082: outdata = 32'd38454;
			27083: outdata = 32'd38453;
			27084: outdata = 32'd38452;
			27085: outdata = 32'd38451;
			27086: outdata = 32'd38450;
			27087: outdata = 32'd38449;
			27088: outdata = 32'd38448;
			27089: outdata = 32'd38447;
			27090: outdata = 32'd38446;
			27091: outdata = 32'd38445;
			27092: outdata = 32'd38444;
			27093: outdata = 32'd38443;
			27094: outdata = 32'd38442;
			27095: outdata = 32'd38441;
			27096: outdata = 32'd38440;
			27097: outdata = 32'd38439;
			27098: outdata = 32'd38438;
			27099: outdata = 32'd38437;
			27100: outdata = 32'd38436;
			27101: outdata = 32'd38435;
			27102: outdata = 32'd38434;
			27103: outdata = 32'd38433;
			27104: outdata = 32'd38432;
			27105: outdata = 32'd38431;
			27106: outdata = 32'd38430;
			27107: outdata = 32'd38429;
			27108: outdata = 32'd38428;
			27109: outdata = 32'd38427;
			27110: outdata = 32'd38426;
			27111: outdata = 32'd38425;
			27112: outdata = 32'd38424;
			27113: outdata = 32'd38423;
			27114: outdata = 32'd38422;
			27115: outdata = 32'd38421;
			27116: outdata = 32'd38420;
			27117: outdata = 32'd38419;
			27118: outdata = 32'd38418;
			27119: outdata = 32'd38417;
			27120: outdata = 32'd38416;
			27121: outdata = 32'd38415;
			27122: outdata = 32'd38414;
			27123: outdata = 32'd38413;
			27124: outdata = 32'd38412;
			27125: outdata = 32'd38411;
			27126: outdata = 32'd38410;
			27127: outdata = 32'd38409;
			27128: outdata = 32'd38408;
			27129: outdata = 32'd38407;
			27130: outdata = 32'd38406;
			27131: outdata = 32'd38405;
			27132: outdata = 32'd38404;
			27133: outdata = 32'd38403;
			27134: outdata = 32'd38402;
			27135: outdata = 32'd38401;
			27136: outdata = 32'd38400;
			27137: outdata = 32'd38399;
			27138: outdata = 32'd38398;
			27139: outdata = 32'd38397;
			27140: outdata = 32'd38396;
			27141: outdata = 32'd38395;
			27142: outdata = 32'd38394;
			27143: outdata = 32'd38393;
			27144: outdata = 32'd38392;
			27145: outdata = 32'd38391;
			27146: outdata = 32'd38390;
			27147: outdata = 32'd38389;
			27148: outdata = 32'd38388;
			27149: outdata = 32'd38387;
			27150: outdata = 32'd38386;
			27151: outdata = 32'd38385;
			27152: outdata = 32'd38384;
			27153: outdata = 32'd38383;
			27154: outdata = 32'd38382;
			27155: outdata = 32'd38381;
			27156: outdata = 32'd38380;
			27157: outdata = 32'd38379;
			27158: outdata = 32'd38378;
			27159: outdata = 32'd38377;
			27160: outdata = 32'd38376;
			27161: outdata = 32'd38375;
			27162: outdata = 32'd38374;
			27163: outdata = 32'd38373;
			27164: outdata = 32'd38372;
			27165: outdata = 32'd38371;
			27166: outdata = 32'd38370;
			27167: outdata = 32'd38369;
			27168: outdata = 32'd38368;
			27169: outdata = 32'd38367;
			27170: outdata = 32'd38366;
			27171: outdata = 32'd38365;
			27172: outdata = 32'd38364;
			27173: outdata = 32'd38363;
			27174: outdata = 32'd38362;
			27175: outdata = 32'd38361;
			27176: outdata = 32'd38360;
			27177: outdata = 32'd38359;
			27178: outdata = 32'd38358;
			27179: outdata = 32'd38357;
			27180: outdata = 32'd38356;
			27181: outdata = 32'd38355;
			27182: outdata = 32'd38354;
			27183: outdata = 32'd38353;
			27184: outdata = 32'd38352;
			27185: outdata = 32'd38351;
			27186: outdata = 32'd38350;
			27187: outdata = 32'd38349;
			27188: outdata = 32'd38348;
			27189: outdata = 32'd38347;
			27190: outdata = 32'd38346;
			27191: outdata = 32'd38345;
			27192: outdata = 32'd38344;
			27193: outdata = 32'd38343;
			27194: outdata = 32'd38342;
			27195: outdata = 32'd38341;
			27196: outdata = 32'd38340;
			27197: outdata = 32'd38339;
			27198: outdata = 32'd38338;
			27199: outdata = 32'd38337;
			27200: outdata = 32'd38336;
			27201: outdata = 32'd38335;
			27202: outdata = 32'd38334;
			27203: outdata = 32'd38333;
			27204: outdata = 32'd38332;
			27205: outdata = 32'd38331;
			27206: outdata = 32'd38330;
			27207: outdata = 32'd38329;
			27208: outdata = 32'd38328;
			27209: outdata = 32'd38327;
			27210: outdata = 32'd38326;
			27211: outdata = 32'd38325;
			27212: outdata = 32'd38324;
			27213: outdata = 32'd38323;
			27214: outdata = 32'd38322;
			27215: outdata = 32'd38321;
			27216: outdata = 32'd38320;
			27217: outdata = 32'd38319;
			27218: outdata = 32'd38318;
			27219: outdata = 32'd38317;
			27220: outdata = 32'd38316;
			27221: outdata = 32'd38315;
			27222: outdata = 32'd38314;
			27223: outdata = 32'd38313;
			27224: outdata = 32'd38312;
			27225: outdata = 32'd38311;
			27226: outdata = 32'd38310;
			27227: outdata = 32'd38309;
			27228: outdata = 32'd38308;
			27229: outdata = 32'd38307;
			27230: outdata = 32'd38306;
			27231: outdata = 32'd38305;
			27232: outdata = 32'd38304;
			27233: outdata = 32'd38303;
			27234: outdata = 32'd38302;
			27235: outdata = 32'd38301;
			27236: outdata = 32'd38300;
			27237: outdata = 32'd38299;
			27238: outdata = 32'd38298;
			27239: outdata = 32'd38297;
			27240: outdata = 32'd38296;
			27241: outdata = 32'd38295;
			27242: outdata = 32'd38294;
			27243: outdata = 32'd38293;
			27244: outdata = 32'd38292;
			27245: outdata = 32'd38291;
			27246: outdata = 32'd38290;
			27247: outdata = 32'd38289;
			27248: outdata = 32'd38288;
			27249: outdata = 32'd38287;
			27250: outdata = 32'd38286;
			27251: outdata = 32'd38285;
			27252: outdata = 32'd38284;
			27253: outdata = 32'd38283;
			27254: outdata = 32'd38282;
			27255: outdata = 32'd38281;
			27256: outdata = 32'd38280;
			27257: outdata = 32'd38279;
			27258: outdata = 32'd38278;
			27259: outdata = 32'd38277;
			27260: outdata = 32'd38276;
			27261: outdata = 32'd38275;
			27262: outdata = 32'd38274;
			27263: outdata = 32'd38273;
			27264: outdata = 32'd38272;
			27265: outdata = 32'd38271;
			27266: outdata = 32'd38270;
			27267: outdata = 32'd38269;
			27268: outdata = 32'd38268;
			27269: outdata = 32'd38267;
			27270: outdata = 32'd38266;
			27271: outdata = 32'd38265;
			27272: outdata = 32'd38264;
			27273: outdata = 32'd38263;
			27274: outdata = 32'd38262;
			27275: outdata = 32'd38261;
			27276: outdata = 32'd38260;
			27277: outdata = 32'd38259;
			27278: outdata = 32'd38258;
			27279: outdata = 32'd38257;
			27280: outdata = 32'd38256;
			27281: outdata = 32'd38255;
			27282: outdata = 32'd38254;
			27283: outdata = 32'd38253;
			27284: outdata = 32'd38252;
			27285: outdata = 32'd38251;
			27286: outdata = 32'd38250;
			27287: outdata = 32'd38249;
			27288: outdata = 32'd38248;
			27289: outdata = 32'd38247;
			27290: outdata = 32'd38246;
			27291: outdata = 32'd38245;
			27292: outdata = 32'd38244;
			27293: outdata = 32'd38243;
			27294: outdata = 32'd38242;
			27295: outdata = 32'd38241;
			27296: outdata = 32'd38240;
			27297: outdata = 32'd38239;
			27298: outdata = 32'd38238;
			27299: outdata = 32'd38237;
			27300: outdata = 32'd38236;
			27301: outdata = 32'd38235;
			27302: outdata = 32'd38234;
			27303: outdata = 32'd38233;
			27304: outdata = 32'd38232;
			27305: outdata = 32'd38231;
			27306: outdata = 32'd38230;
			27307: outdata = 32'd38229;
			27308: outdata = 32'd38228;
			27309: outdata = 32'd38227;
			27310: outdata = 32'd38226;
			27311: outdata = 32'd38225;
			27312: outdata = 32'd38224;
			27313: outdata = 32'd38223;
			27314: outdata = 32'd38222;
			27315: outdata = 32'd38221;
			27316: outdata = 32'd38220;
			27317: outdata = 32'd38219;
			27318: outdata = 32'd38218;
			27319: outdata = 32'd38217;
			27320: outdata = 32'd38216;
			27321: outdata = 32'd38215;
			27322: outdata = 32'd38214;
			27323: outdata = 32'd38213;
			27324: outdata = 32'd38212;
			27325: outdata = 32'd38211;
			27326: outdata = 32'd38210;
			27327: outdata = 32'd38209;
			27328: outdata = 32'd38208;
			27329: outdata = 32'd38207;
			27330: outdata = 32'd38206;
			27331: outdata = 32'd38205;
			27332: outdata = 32'd38204;
			27333: outdata = 32'd38203;
			27334: outdata = 32'd38202;
			27335: outdata = 32'd38201;
			27336: outdata = 32'd38200;
			27337: outdata = 32'd38199;
			27338: outdata = 32'd38198;
			27339: outdata = 32'd38197;
			27340: outdata = 32'd38196;
			27341: outdata = 32'd38195;
			27342: outdata = 32'd38194;
			27343: outdata = 32'd38193;
			27344: outdata = 32'd38192;
			27345: outdata = 32'd38191;
			27346: outdata = 32'd38190;
			27347: outdata = 32'd38189;
			27348: outdata = 32'd38188;
			27349: outdata = 32'd38187;
			27350: outdata = 32'd38186;
			27351: outdata = 32'd38185;
			27352: outdata = 32'd38184;
			27353: outdata = 32'd38183;
			27354: outdata = 32'd38182;
			27355: outdata = 32'd38181;
			27356: outdata = 32'd38180;
			27357: outdata = 32'd38179;
			27358: outdata = 32'd38178;
			27359: outdata = 32'd38177;
			27360: outdata = 32'd38176;
			27361: outdata = 32'd38175;
			27362: outdata = 32'd38174;
			27363: outdata = 32'd38173;
			27364: outdata = 32'd38172;
			27365: outdata = 32'd38171;
			27366: outdata = 32'd38170;
			27367: outdata = 32'd38169;
			27368: outdata = 32'd38168;
			27369: outdata = 32'd38167;
			27370: outdata = 32'd38166;
			27371: outdata = 32'd38165;
			27372: outdata = 32'd38164;
			27373: outdata = 32'd38163;
			27374: outdata = 32'd38162;
			27375: outdata = 32'd38161;
			27376: outdata = 32'd38160;
			27377: outdata = 32'd38159;
			27378: outdata = 32'd38158;
			27379: outdata = 32'd38157;
			27380: outdata = 32'd38156;
			27381: outdata = 32'd38155;
			27382: outdata = 32'd38154;
			27383: outdata = 32'd38153;
			27384: outdata = 32'd38152;
			27385: outdata = 32'd38151;
			27386: outdata = 32'd38150;
			27387: outdata = 32'd38149;
			27388: outdata = 32'd38148;
			27389: outdata = 32'd38147;
			27390: outdata = 32'd38146;
			27391: outdata = 32'd38145;
			27392: outdata = 32'd38144;
			27393: outdata = 32'd38143;
			27394: outdata = 32'd38142;
			27395: outdata = 32'd38141;
			27396: outdata = 32'd38140;
			27397: outdata = 32'd38139;
			27398: outdata = 32'd38138;
			27399: outdata = 32'd38137;
			27400: outdata = 32'd38136;
			27401: outdata = 32'd38135;
			27402: outdata = 32'd38134;
			27403: outdata = 32'd38133;
			27404: outdata = 32'd38132;
			27405: outdata = 32'd38131;
			27406: outdata = 32'd38130;
			27407: outdata = 32'd38129;
			27408: outdata = 32'd38128;
			27409: outdata = 32'd38127;
			27410: outdata = 32'd38126;
			27411: outdata = 32'd38125;
			27412: outdata = 32'd38124;
			27413: outdata = 32'd38123;
			27414: outdata = 32'd38122;
			27415: outdata = 32'd38121;
			27416: outdata = 32'd38120;
			27417: outdata = 32'd38119;
			27418: outdata = 32'd38118;
			27419: outdata = 32'd38117;
			27420: outdata = 32'd38116;
			27421: outdata = 32'd38115;
			27422: outdata = 32'd38114;
			27423: outdata = 32'd38113;
			27424: outdata = 32'd38112;
			27425: outdata = 32'd38111;
			27426: outdata = 32'd38110;
			27427: outdata = 32'd38109;
			27428: outdata = 32'd38108;
			27429: outdata = 32'd38107;
			27430: outdata = 32'd38106;
			27431: outdata = 32'd38105;
			27432: outdata = 32'd38104;
			27433: outdata = 32'd38103;
			27434: outdata = 32'd38102;
			27435: outdata = 32'd38101;
			27436: outdata = 32'd38100;
			27437: outdata = 32'd38099;
			27438: outdata = 32'd38098;
			27439: outdata = 32'd38097;
			27440: outdata = 32'd38096;
			27441: outdata = 32'd38095;
			27442: outdata = 32'd38094;
			27443: outdata = 32'd38093;
			27444: outdata = 32'd38092;
			27445: outdata = 32'd38091;
			27446: outdata = 32'd38090;
			27447: outdata = 32'd38089;
			27448: outdata = 32'd38088;
			27449: outdata = 32'd38087;
			27450: outdata = 32'd38086;
			27451: outdata = 32'd38085;
			27452: outdata = 32'd38084;
			27453: outdata = 32'd38083;
			27454: outdata = 32'd38082;
			27455: outdata = 32'd38081;
			27456: outdata = 32'd38080;
			27457: outdata = 32'd38079;
			27458: outdata = 32'd38078;
			27459: outdata = 32'd38077;
			27460: outdata = 32'd38076;
			27461: outdata = 32'd38075;
			27462: outdata = 32'd38074;
			27463: outdata = 32'd38073;
			27464: outdata = 32'd38072;
			27465: outdata = 32'd38071;
			27466: outdata = 32'd38070;
			27467: outdata = 32'd38069;
			27468: outdata = 32'd38068;
			27469: outdata = 32'd38067;
			27470: outdata = 32'd38066;
			27471: outdata = 32'd38065;
			27472: outdata = 32'd38064;
			27473: outdata = 32'd38063;
			27474: outdata = 32'd38062;
			27475: outdata = 32'd38061;
			27476: outdata = 32'd38060;
			27477: outdata = 32'd38059;
			27478: outdata = 32'd38058;
			27479: outdata = 32'd38057;
			27480: outdata = 32'd38056;
			27481: outdata = 32'd38055;
			27482: outdata = 32'd38054;
			27483: outdata = 32'd38053;
			27484: outdata = 32'd38052;
			27485: outdata = 32'd38051;
			27486: outdata = 32'd38050;
			27487: outdata = 32'd38049;
			27488: outdata = 32'd38048;
			27489: outdata = 32'd38047;
			27490: outdata = 32'd38046;
			27491: outdata = 32'd38045;
			27492: outdata = 32'd38044;
			27493: outdata = 32'd38043;
			27494: outdata = 32'd38042;
			27495: outdata = 32'd38041;
			27496: outdata = 32'd38040;
			27497: outdata = 32'd38039;
			27498: outdata = 32'd38038;
			27499: outdata = 32'd38037;
			27500: outdata = 32'd38036;
			27501: outdata = 32'd38035;
			27502: outdata = 32'd38034;
			27503: outdata = 32'd38033;
			27504: outdata = 32'd38032;
			27505: outdata = 32'd38031;
			27506: outdata = 32'd38030;
			27507: outdata = 32'd38029;
			27508: outdata = 32'd38028;
			27509: outdata = 32'd38027;
			27510: outdata = 32'd38026;
			27511: outdata = 32'd38025;
			27512: outdata = 32'd38024;
			27513: outdata = 32'd38023;
			27514: outdata = 32'd38022;
			27515: outdata = 32'd38021;
			27516: outdata = 32'd38020;
			27517: outdata = 32'd38019;
			27518: outdata = 32'd38018;
			27519: outdata = 32'd38017;
			27520: outdata = 32'd38016;
			27521: outdata = 32'd38015;
			27522: outdata = 32'd38014;
			27523: outdata = 32'd38013;
			27524: outdata = 32'd38012;
			27525: outdata = 32'd38011;
			27526: outdata = 32'd38010;
			27527: outdata = 32'd38009;
			27528: outdata = 32'd38008;
			27529: outdata = 32'd38007;
			27530: outdata = 32'd38006;
			27531: outdata = 32'd38005;
			27532: outdata = 32'd38004;
			27533: outdata = 32'd38003;
			27534: outdata = 32'd38002;
			27535: outdata = 32'd38001;
			27536: outdata = 32'd38000;
			27537: outdata = 32'd37999;
			27538: outdata = 32'd37998;
			27539: outdata = 32'd37997;
			27540: outdata = 32'd37996;
			27541: outdata = 32'd37995;
			27542: outdata = 32'd37994;
			27543: outdata = 32'd37993;
			27544: outdata = 32'd37992;
			27545: outdata = 32'd37991;
			27546: outdata = 32'd37990;
			27547: outdata = 32'd37989;
			27548: outdata = 32'd37988;
			27549: outdata = 32'd37987;
			27550: outdata = 32'd37986;
			27551: outdata = 32'd37985;
			27552: outdata = 32'd37984;
			27553: outdata = 32'd37983;
			27554: outdata = 32'd37982;
			27555: outdata = 32'd37981;
			27556: outdata = 32'd37980;
			27557: outdata = 32'd37979;
			27558: outdata = 32'd37978;
			27559: outdata = 32'd37977;
			27560: outdata = 32'd37976;
			27561: outdata = 32'd37975;
			27562: outdata = 32'd37974;
			27563: outdata = 32'd37973;
			27564: outdata = 32'd37972;
			27565: outdata = 32'd37971;
			27566: outdata = 32'd37970;
			27567: outdata = 32'd37969;
			27568: outdata = 32'd37968;
			27569: outdata = 32'd37967;
			27570: outdata = 32'd37966;
			27571: outdata = 32'd37965;
			27572: outdata = 32'd37964;
			27573: outdata = 32'd37963;
			27574: outdata = 32'd37962;
			27575: outdata = 32'd37961;
			27576: outdata = 32'd37960;
			27577: outdata = 32'd37959;
			27578: outdata = 32'd37958;
			27579: outdata = 32'd37957;
			27580: outdata = 32'd37956;
			27581: outdata = 32'd37955;
			27582: outdata = 32'd37954;
			27583: outdata = 32'd37953;
			27584: outdata = 32'd37952;
			27585: outdata = 32'd37951;
			27586: outdata = 32'd37950;
			27587: outdata = 32'd37949;
			27588: outdata = 32'd37948;
			27589: outdata = 32'd37947;
			27590: outdata = 32'd37946;
			27591: outdata = 32'd37945;
			27592: outdata = 32'd37944;
			27593: outdata = 32'd37943;
			27594: outdata = 32'd37942;
			27595: outdata = 32'd37941;
			27596: outdata = 32'd37940;
			27597: outdata = 32'd37939;
			27598: outdata = 32'd37938;
			27599: outdata = 32'd37937;
			27600: outdata = 32'd37936;
			27601: outdata = 32'd37935;
			27602: outdata = 32'd37934;
			27603: outdata = 32'd37933;
			27604: outdata = 32'd37932;
			27605: outdata = 32'd37931;
			27606: outdata = 32'd37930;
			27607: outdata = 32'd37929;
			27608: outdata = 32'd37928;
			27609: outdata = 32'd37927;
			27610: outdata = 32'd37926;
			27611: outdata = 32'd37925;
			27612: outdata = 32'd37924;
			27613: outdata = 32'd37923;
			27614: outdata = 32'd37922;
			27615: outdata = 32'd37921;
			27616: outdata = 32'd37920;
			27617: outdata = 32'd37919;
			27618: outdata = 32'd37918;
			27619: outdata = 32'd37917;
			27620: outdata = 32'd37916;
			27621: outdata = 32'd37915;
			27622: outdata = 32'd37914;
			27623: outdata = 32'd37913;
			27624: outdata = 32'd37912;
			27625: outdata = 32'd37911;
			27626: outdata = 32'd37910;
			27627: outdata = 32'd37909;
			27628: outdata = 32'd37908;
			27629: outdata = 32'd37907;
			27630: outdata = 32'd37906;
			27631: outdata = 32'd37905;
			27632: outdata = 32'd37904;
			27633: outdata = 32'd37903;
			27634: outdata = 32'd37902;
			27635: outdata = 32'd37901;
			27636: outdata = 32'd37900;
			27637: outdata = 32'd37899;
			27638: outdata = 32'd37898;
			27639: outdata = 32'd37897;
			27640: outdata = 32'd37896;
			27641: outdata = 32'd37895;
			27642: outdata = 32'd37894;
			27643: outdata = 32'd37893;
			27644: outdata = 32'd37892;
			27645: outdata = 32'd37891;
			27646: outdata = 32'd37890;
			27647: outdata = 32'd37889;
			27648: outdata = 32'd37888;
			27649: outdata = 32'd37887;
			27650: outdata = 32'd37886;
			27651: outdata = 32'd37885;
			27652: outdata = 32'd37884;
			27653: outdata = 32'd37883;
			27654: outdata = 32'd37882;
			27655: outdata = 32'd37881;
			27656: outdata = 32'd37880;
			27657: outdata = 32'd37879;
			27658: outdata = 32'd37878;
			27659: outdata = 32'd37877;
			27660: outdata = 32'd37876;
			27661: outdata = 32'd37875;
			27662: outdata = 32'd37874;
			27663: outdata = 32'd37873;
			27664: outdata = 32'd37872;
			27665: outdata = 32'd37871;
			27666: outdata = 32'd37870;
			27667: outdata = 32'd37869;
			27668: outdata = 32'd37868;
			27669: outdata = 32'd37867;
			27670: outdata = 32'd37866;
			27671: outdata = 32'd37865;
			27672: outdata = 32'd37864;
			27673: outdata = 32'd37863;
			27674: outdata = 32'd37862;
			27675: outdata = 32'd37861;
			27676: outdata = 32'd37860;
			27677: outdata = 32'd37859;
			27678: outdata = 32'd37858;
			27679: outdata = 32'd37857;
			27680: outdata = 32'd37856;
			27681: outdata = 32'd37855;
			27682: outdata = 32'd37854;
			27683: outdata = 32'd37853;
			27684: outdata = 32'd37852;
			27685: outdata = 32'd37851;
			27686: outdata = 32'd37850;
			27687: outdata = 32'd37849;
			27688: outdata = 32'd37848;
			27689: outdata = 32'd37847;
			27690: outdata = 32'd37846;
			27691: outdata = 32'd37845;
			27692: outdata = 32'd37844;
			27693: outdata = 32'd37843;
			27694: outdata = 32'd37842;
			27695: outdata = 32'd37841;
			27696: outdata = 32'd37840;
			27697: outdata = 32'd37839;
			27698: outdata = 32'd37838;
			27699: outdata = 32'd37837;
			27700: outdata = 32'd37836;
			27701: outdata = 32'd37835;
			27702: outdata = 32'd37834;
			27703: outdata = 32'd37833;
			27704: outdata = 32'd37832;
			27705: outdata = 32'd37831;
			27706: outdata = 32'd37830;
			27707: outdata = 32'd37829;
			27708: outdata = 32'd37828;
			27709: outdata = 32'd37827;
			27710: outdata = 32'd37826;
			27711: outdata = 32'd37825;
			27712: outdata = 32'd37824;
			27713: outdata = 32'd37823;
			27714: outdata = 32'd37822;
			27715: outdata = 32'd37821;
			27716: outdata = 32'd37820;
			27717: outdata = 32'd37819;
			27718: outdata = 32'd37818;
			27719: outdata = 32'd37817;
			27720: outdata = 32'd37816;
			27721: outdata = 32'd37815;
			27722: outdata = 32'd37814;
			27723: outdata = 32'd37813;
			27724: outdata = 32'd37812;
			27725: outdata = 32'd37811;
			27726: outdata = 32'd37810;
			27727: outdata = 32'd37809;
			27728: outdata = 32'd37808;
			27729: outdata = 32'd37807;
			27730: outdata = 32'd37806;
			27731: outdata = 32'd37805;
			27732: outdata = 32'd37804;
			27733: outdata = 32'd37803;
			27734: outdata = 32'd37802;
			27735: outdata = 32'd37801;
			27736: outdata = 32'd37800;
			27737: outdata = 32'd37799;
			27738: outdata = 32'd37798;
			27739: outdata = 32'd37797;
			27740: outdata = 32'd37796;
			27741: outdata = 32'd37795;
			27742: outdata = 32'd37794;
			27743: outdata = 32'd37793;
			27744: outdata = 32'd37792;
			27745: outdata = 32'd37791;
			27746: outdata = 32'd37790;
			27747: outdata = 32'd37789;
			27748: outdata = 32'd37788;
			27749: outdata = 32'd37787;
			27750: outdata = 32'd37786;
			27751: outdata = 32'd37785;
			27752: outdata = 32'd37784;
			27753: outdata = 32'd37783;
			27754: outdata = 32'd37782;
			27755: outdata = 32'd37781;
			27756: outdata = 32'd37780;
			27757: outdata = 32'd37779;
			27758: outdata = 32'd37778;
			27759: outdata = 32'd37777;
			27760: outdata = 32'd37776;
			27761: outdata = 32'd37775;
			27762: outdata = 32'd37774;
			27763: outdata = 32'd37773;
			27764: outdata = 32'd37772;
			27765: outdata = 32'd37771;
			27766: outdata = 32'd37770;
			27767: outdata = 32'd37769;
			27768: outdata = 32'd37768;
			27769: outdata = 32'd37767;
			27770: outdata = 32'd37766;
			27771: outdata = 32'd37765;
			27772: outdata = 32'd37764;
			27773: outdata = 32'd37763;
			27774: outdata = 32'd37762;
			27775: outdata = 32'd37761;
			27776: outdata = 32'd37760;
			27777: outdata = 32'd37759;
			27778: outdata = 32'd37758;
			27779: outdata = 32'd37757;
			27780: outdata = 32'd37756;
			27781: outdata = 32'd37755;
			27782: outdata = 32'd37754;
			27783: outdata = 32'd37753;
			27784: outdata = 32'd37752;
			27785: outdata = 32'd37751;
			27786: outdata = 32'd37750;
			27787: outdata = 32'd37749;
			27788: outdata = 32'd37748;
			27789: outdata = 32'd37747;
			27790: outdata = 32'd37746;
			27791: outdata = 32'd37745;
			27792: outdata = 32'd37744;
			27793: outdata = 32'd37743;
			27794: outdata = 32'd37742;
			27795: outdata = 32'd37741;
			27796: outdata = 32'd37740;
			27797: outdata = 32'd37739;
			27798: outdata = 32'd37738;
			27799: outdata = 32'd37737;
			27800: outdata = 32'd37736;
			27801: outdata = 32'd37735;
			27802: outdata = 32'd37734;
			27803: outdata = 32'd37733;
			27804: outdata = 32'd37732;
			27805: outdata = 32'd37731;
			27806: outdata = 32'd37730;
			27807: outdata = 32'd37729;
			27808: outdata = 32'd37728;
			27809: outdata = 32'd37727;
			27810: outdata = 32'd37726;
			27811: outdata = 32'd37725;
			27812: outdata = 32'd37724;
			27813: outdata = 32'd37723;
			27814: outdata = 32'd37722;
			27815: outdata = 32'd37721;
			27816: outdata = 32'd37720;
			27817: outdata = 32'd37719;
			27818: outdata = 32'd37718;
			27819: outdata = 32'd37717;
			27820: outdata = 32'd37716;
			27821: outdata = 32'd37715;
			27822: outdata = 32'd37714;
			27823: outdata = 32'd37713;
			27824: outdata = 32'd37712;
			27825: outdata = 32'd37711;
			27826: outdata = 32'd37710;
			27827: outdata = 32'd37709;
			27828: outdata = 32'd37708;
			27829: outdata = 32'd37707;
			27830: outdata = 32'd37706;
			27831: outdata = 32'd37705;
			27832: outdata = 32'd37704;
			27833: outdata = 32'd37703;
			27834: outdata = 32'd37702;
			27835: outdata = 32'd37701;
			27836: outdata = 32'd37700;
			27837: outdata = 32'd37699;
			27838: outdata = 32'd37698;
			27839: outdata = 32'd37697;
			27840: outdata = 32'd37696;
			27841: outdata = 32'd37695;
			27842: outdata = 32'd37694;
			27843: outdata = 32'd37693;
			27844: outdata = 32'd37692;
			27845: outdata = 32'd37691;
			27846: outdata = 32'd37690;
			27847: outdata = 32'd37689;
			27848: outdata = 32'd37688;
			27849: outdata = 32'd37687;
			27850: outdata = 32'd37686;
			27851: outdata = 32'd37685;
			27852: outdata = 32'd37684;
			27853: outdata = 32'd37683;
			27854: outdata = 32'd37682;
			27855: outdata = 32'd37681;
			27856: outdata = 32'd37680;
			27857: outdata = 32'd37679;
			27858: outdata = 32'd37678;
			27859: outdata = 32'd37677;
			27860: outdata = 32'd37676;
			27861: outdata = 32'd37675;
			27862: outdata = 32'd37674;
			27863: outdata = 32'd37673;
			27864: outdata = 32'd37672;
			27865: outdata = 32'd37671;
			27866: outdata = 32'd37670;
			27867: outdata = 32'd37669;
			27868: outdata = 32'd37668;
			27869: outdata = 32'd37667;
			27870: outdata = 32'd37666;
			27871: outdata = 32'd37665;
			27872: outdata = 32'd37664;
			27873: outdata = 32'd37663;
			27874: outdata = 32'd37662;
			27875: outdata = 32'd37661;
			27876: outdata = 32'd37660;
			27877: outdata = 32'd37659;
			27878: outdata = 32'd37658;
			27879: outdata = 32'd37657;
			27880: outdata = 32'd37656;
			27881: outdata = 32'd37655;
			27882: outdata = 32'd37654;
			27883: outdata = 32'd37653;
			27884: outdata = 32'd37652;
			27885: outdata = 32'd37651;
			27886: outdata = 32'd37650;
			27887: outdata = 32'd37649;
			27888: outdata = 32'd37648;
			27889: outdata = 32'd37647;
			27890: outdata = 32'd37646;
			27891: outdata = 32'd37645;
			27892: outdata = 32'd37644;
			27893: outdata = 32'd37643;
			27894: outdata = 32'd37642;
			27895: outdata = 32'd37641;
			27896: outdata = 32'd37640;
			27897: outdata = 32'd37639;
			27898: outdata = 32'd37638;
			27899: outdata = 32'd37637;
			27900: outdata = 32'd37636;
			27901: outdata = 32'd37635;
			27902: outdata = 32'd37634;
			27903: outdata = 32'd37633;
			27904: outdata = 32'd37632;
			27905: outdata = 32'd37631;
			27906: outdata = 32'd37630;
			27907: outdata = 32'd37629;
			27908: outdata = 32'd37628;
			27909: outdata = 32'd37627;
			27910: outdata = 32'd37626;
			27911: outdata = 32'd37625;
			27912: outdata = 32'd37624;
			27913: outdata = 32'd37623;
			27914: outdata = 32'd37622;
			27915: outdata = 32'd37621;
			27916: outdata = 32'd37620;
			27917: outdata = 32'd37619;
			27918: outdata = 32'd37618;
			27919: outdata = 32'd37617;
			27920: outdata = 32'd37616;
			27921: outdata = 32'd37615;
			27922: outdata = 32'd37614;
			27923: outdata = 32'd37613;
			27924: outdata = 32'd37612;
			27925: outdata = 32'd37611;
			27926: outdata = 32'd37610;
			27927: outdata = 32'd37609;
			27928: outdata = 32'd37608;
			27929: outdata = 32'd37607;
			27930: outdata = 32'd37606;
			27931: outdata = 32'd37605;
			27932: outdata = 32'd37604;
			27933: outdata = 32'd37603;
			27934: outdata = 32'd37602;
			27935: outdata = 32'd37601;
			27936: outdata = 32'd37600;
			27937: outdata = 32'd37599;
			27938: outdata = 32'd37598;
			27939: outdata = 32'd37597;
			27940: outdata = 32'd37596;
			27941: outdata = 32'd37595;
			27942: outdata = 32'd37594;
			27943: outdata = 32'd37593;
			27944: outdata = 32'd37592;
			27945: outdata = 32'd37591;
			27946: outdata = 32'd37590;
			27947: outdata = 32'd37589;
			27948: outdata = 32'd37588;
			27949: outdata = 32'd37587;
			27950: outdata = 32'd37586;
			27951: outdata = 32'd37585;
			27952: outdata = 32'd37584;
			27953: outdata = 32'd37583;
			27954: outdata = 32'd37582;
			27955: outdata = 32'd37581;
			27956: outdata = 32'd37580;
			27957: outdata = 32'd37579;
			27958: outdata = 32'd37578;
			27959: outdata = 32'd37577;
			27960: outdata = 32'd37576;
			27961: outdata = 32'd37575;
			27962: outdata = 32'd37574;
			27963: outdata = 32'd37573;
			27964: outdata = 32'd37572;
			27965: outdata = 32'd37571;
			27966: outdata = 32'd37570;
			27967: outdata = 32'd37569;
			27968: outdata = 32'd37568;
			27969: outdata = 32'd37567;
			27970: outdata = 32'd37566;
			27971: outdata = 32'd37565;
			27972: outdata = 32'd37564;
			27973: outdata = 32'd37563;
			27974: outdata = 32'd37562;
			27975: outdata = 32'd37561;
			27976: outdata = 32'd37560;
			27977: outdata = 32'd37559;
			27978: outdata = 32'd37558;
			27979: outdata = 32'd37557;
			27980: outdata = 32'd37556;
			27981: outdata = 32'd37555;
			27982: outdata = 32'd37554;
			27983: outdata = 32'd37553;
			27984: outdata = 32'd37552;
			27985: outdata = 32'd37551;
			27986: outdata = 32'd37550;
			27987: outdata = 32'd37549;
			27988: outdata = 32'd37548;
			27989: outdata = 32'd37547;
			27990: outdata = 32'd37546;
			27991: outdata = 32'd37545;
			27992: outdata = 32'd37544;
			27993: outdata = 32'd37543;
			27994: outdata = 32'd37542;
			27995: outdata = 32'd37541;
			27996: outdata = 32'd37540;
			27997: outdata = 32'd37539;
			27998: outdata = 32'd37538;
			27999: outdata = 32'd37537;
			28000: outdata = 32'd37536;
			28001: outdata = 32'd37535;
			28002: outdata = 32'd37534;
			28003: outdata = 32'd37533;
			28004: outdata = 32'd37532;
			28005: outdata = 32'd37531;
			28006: outdata = 32'd37530;
			28007: outdata = 32'd37529;
			28008: outdata = 32'd37528;
			28009: outdata = 32'd37527;
			28010: outdata = 32'd37526;
			28011: outdata = 32'd37525;
			28012: outdata = 32'd37524;
			28013: outdata = 32'd37523;
			28014: outdata = 32'd37522;
			28015: outdata = 32'd37521;
			28016: outdata = 32'd37520;
			28017: outdata = 32'd37519;
			28018: outdata = 32'd37518;
			28019: outdata = 32'd37517;
			28020: outdata = 32'd37516;
			28021: outdata = 32'd37515;
			28022: outdata = 32'd37514;
			28023: outdata = 32'd37513;
			28024: outdata = 32'd37512;
			28025: outdata = 32'd37511;
			28026: outdata = 32'd37510;
			28027: outdata = 32'd37509;
			28028: outdata = 32'd37508;
			28029: outdata = 32'd37507;
			28030: outdata = 32'd37506;
			28031: outdata = 32'd37505;
			28032: outdata = 32'd37504;
			28033: outdata = 32'd37503;
			28034: outdata = 32'd37502;
			28035: outdata = 32'd37501;
			28036: outdata = 32'd37500;
			28037: outdata = 32'd37499;
			28038: outdata = 32'd37498;
			28039: outdata = 32'd37497;
			28040: outdata = 32'd37496;
			28041: outdata = 32'd37495;
			28042: outdata = 32'd37494;
			28043: outdata = 32'd37493;
			28044: outdata = 32'd37492;
			28045: outdata = 32'd37491;
			28046: outdata = 32'd37490;
			28047: outdata = 32'd37489;
			28048: outdata = 32'd37488;
			28049: outdata = 32'd37487;
			28050: outdata = 32'd37486;
			28051: outdata = 32'd37485;
			28052: outdata = 32'd37484;
			28053: outdata = 32'd37483;
			28054: outdata = 32'd37482;
			28055: outdata = 32'd37481;
			28056: outdata = 32'd37480;
			28057: outdata = 32'd37479;
			28058: outdata = 32'd37478;
			28059: outdata = 32'd37477;
			28060: outdata = 32'd37476;
			28061: outdata = 32'd37475;
			28062: outdata = 32'd37474;
			28063: outdata = 32'd37473;
			28064: outdata = 32'd37472;
			28065: outdata = 32'd37471;
			28066: outdata = 32'd37470;
			28067: outdata = 32'd37469;
			28068: outdata = 32'd37468;
			28069: outdata = 32'd37467;
			28070: outdata = 32'd37466;
			28071: outdata = 32'd37465;
			28072: outdata = 32'd37464;
			28073: outdata = 32'd37463;
			28074: outdata = 32'd37462;
			28075: outdata = 32'd37461;
			28076: outdata = 32'd37460;
			28077: outdata = 32'd37459;
			28078: outdata = 32'd37458;
			28079: outdata = 32'd37457;
			28080: outdata = 32'd37456;
			28081: outdata = 32'd37455;
			28082: outdata = 32'd37454;
			28083: outdata = 32'd37453;
			28084: outdata = 32'd37452;
			28085: outdata = 32'd37451;
			28086: outdata = 32'd37450;
			28087: outdata = 32'd37449;
			28088: outdata = 32'd37448;
			28089: outdata = 32'd37447;
			28090: outdata = 32'd37446;
			28091: outdata = 32'd37445;
			28092: outdata = 32'd37444;
			28093: outdata = 32'd37443;
			28094: outdata = 32'd37442;
			28095: outdata = 32'd37441;
			28096: outdata = 32'd37440;
			28097: outdata = 32'd37439;
			28098: outdata = 32'd37438;
			28099: outdata = 32'd37437;
			28100: outdata = 32'd37436;
			28101: outdata = 32'd37435;
			28102: outdata = 32'd37434;
			28103: outdata = 32'd37433;
			28104: outdata = 32'd37432;
			28105: outdata = 32'd37431;
			28106: outdata = 32'd37430;
			28107: outdata = 32'd37429;
			28108: outdata = 32'd37428;
			28109: outdata = 32'd37427;
			28110: outdata = 32'd37426;
			28111: outdata = 32'd37425;
			28112: outdata = 32'd37424;
			28113: outdata = 32'd37423;
			28114: outdata = 32'd37422;
			28115: outdata = 32'd37421;
			28116: outdata = 32'd37420;
			28117: outdata = 32'd37419;
			28118: outdata = 32'd37418;
			28119: outdata = 32'd37417;
			28120: outdata = 32'd37416;
			28121: outdata = 32'd37415;
			28122: outdata = 32'd37414;
			28123: outdata = 32'd37413;
			28124: outdata = 32'd37412;
			28125: outdata = 32'd37411;
			28126: outdata = 32'd37410;
			28127: outdata = 32'd37409;
			28128: outdata = 32'd37408;
			28129: outdata = 32'd37407;
			28130: outdata = 32'd37406;
			28131: outdata = 32'd37405;
			28132: outdata = 32'd37404;
			28133: outdata = 32'd37403;
			28134: outdata = 32'd37402;
			28135: outdata = 32'd37401;
			28136: outdata = 32'd37400;
			28137: outdata = 32'd37399;
			28138: outdata = 32'd37398;
			28139: outdata = 32'd37397;
			28140: outdata = 32'd37396;
			28141: outdata = 32'd37395;
			28142: outdata = 32'd37394;
			28143: outdata = 32'd37393;
			28144: outdata = 32'd37392;
			28145: outdata = 32'd37391;
			28146: outdata = 32'd37390;
			28147: outdata = 32'd37389;
			28148: outdata = 32'd37388;
			28149: outdata = 32'd37387;
			28150: outdata = 32'd37386;
			28151: outdata = 32'd37385;
			28152: outdata = 32'd37384;
			28153: outdata = 32'd37383;
			28154: outdata = 32'd37382;
			28155: outdata = 32'd37381;
			28156: outdata = 32'd37380;
			28157: outdata = 32'd37379;
			28158: outdata = 32'd37378;
			28159: outdata = 32'd37377;
			28160: outdata = 32'd37376;
			28161: outdata = 32'd37375;
			28162: outdata = 32'd37374;
			28163: outdata = 32'd37373;
			28164: outdata = 32'd37372;
			28165: outdata = 32'd37371;
			28166: outdata = 32'd37370;
			28167: outdata = 32'd37369;
			28168: outdata = 32'd37368;
			28169: outdata = 32'd37367;
			28170: outdata = 32'd37366;
			28171: outdata = 32'd37365;
			28172: outdata = 32'd37364;
			28173: outdata = 32'd37363;
			28174: outdata = 32'd37362;
			28175: outdata = 32'd37361;
			28176: outdata = 32'd37360;
			28177: outdata = 32'd37359;
			28178: outdata = 32'd37358;
			28179: outdata = 32'd37357;
			28180: outdata = 32'd37356;
			28181: outdata = 32'd37355;
			28182: outdata = 32'd37354;
			28183: outdata = 32'd37353;
			28184: outdata = 32'd37352;
			28185: outdata = 32'd37351;
			28186: outdata = 32'd37350;
			28187: outdata = 32'd37349;
			28188: outdata = 32'd37348;
			28189: outdata = 32'd37347;
			28190: outdata = 32'd37346;
			28191: outdata = 32'd37345;
			28192: outdata = 32'd37344;
			28193: outdata = 32'd37343;
			28194: outdata = 32'd37342;
			28195: outdata = 32'd37341;
			28196: outdata = 32'd37340;
			28197: outdata = 32'd37339;
			28198: outdata = 32'd37338;
			28199: outdata = 32'd37337;
			28200: outdata = 32'd37336;
			28201: outdata = 32'd37335;
			28202: outdata = 32'd37334;
			28203: outdata = 32'd37333;
			28204: outdata = 32'd37332;
			28205: outdata = 32'd37331;
			28206: outdata = 32'd37330;
			28207: outdata = 32'd37329;
			28208: outdata = 32'd37328;
			28209: outdata = 32'd37327;
			28210: outdata = 32'd37326;
			28211: outdata = 32'd37325;
			28212: outdata = 32'd37324;
			28213: outdata = 32'd37323;
			28214: outdata = 32'd37322;
			28215: outdata = 32'd37321;
			28216: outdata = 32'd37320;
			28217: outdata = 32'd37319;
			28218: outdata = 32'd37318;
			28219: outdata = 32'd37317;
			28220: outdata = 32'd37316;
			28221: outdata = 32'd37315;
			28222: outdata = 32'd37314;
			28223: outdata = 32'd37313;
			28224: outdata = 32'd37312;
			28225: outdata = 32'd37311;
			28226: outdata = 32'd37310;
			28227: outdata = 32'd37309;
			28228: outdata = 32'd37308;
			28229: outdata = 32'd37307;
			28230: outdata = 32'd37306;
			28231: outdata = 32'd37305;
			28232: outdata = 32'd37304;
			28233: outdata = 32'd37303;
			28234: outdata = 32'd37302;
			28235: outdata = 32'd37301;
			28236: outdata = 32'd37300;
			28237: outdata = 32'd37299;
			28238: outdata = 32'd37298;
			28239: outdata = 32'd37297;
			28240: outdata = 32'd37296;
			28241: outdata = 32'd37295;
			28242: outdata = 32'd37294;
			28243: outdata = 32'd37293;
			28244: outdata = 32'd37292;
			28245: outdata = 32'd37291;
			28246: outdata = 32'd37290;
			28247: outdata = 32'd37289;
			28248: outdata = 32'd37288;
			28249: outdata = 32'd37287;
			28250: outdata = 32'd37286;
			28251: outdata = 32'd37285;
			28252: outdata = 32'd37284;
			28253: outdata = 32'd37283;
			28254: outdata = 32'd37282;
			28255: outdata = 32'd37281;
			28256: outdata = 32'd37280;
			28257: outdata = 32'd37279;
			28258: outdata = 32'd37278;
			28259: outdata = 32'd37277;
			28260: outdata = 32'd37276;
			28261: outdata = 32'd37275;
			28262: outdata = 32'd37274;
			28263: outdata = 32'd37273;
			28264: outdata = 32'd37272;
			28265: outdata = 32'd37271;
			28266: outdata = 32'd37270;
			28267: outdata = 32'd37269;
			28268: outdata = 32'd37268;
			28269: outdata = 32'd37267;
			28270: outdata = 32'd37266;
			28271: outdata = 32'd37265;
			28272: outdata = 32'd37264;
			28273: outdata = 32'd37263;
			28274: outdata = 32'd37262;
			28275: outdata = 32'd37261;
			28276: outdata = 32'd37260;
			28277: outdata = 32'd37259;
			28278: outdata = 32'd37258;
			28279: outdata = 32'd37257;
			28280: outdata = 32'd37256;
			28281: outdata = 32'd37255;
			28282: outdata = 32'd37254;
			28283: outdata = 32'd37253;
			28284: outdata = 32'd37252;
			28285: outdata = 32'd37251;
			28286: outdata = 32'd37250;
			28287: outdata = 32'd37249;
			28288: outdata = 32'd37248;
			28289: outdata = 32'd37247;
			28290: outdata = 32'd37246;
			28291: outdata = 32'd37245;
			28292: outdata = 32'd37244;
			28293: outdata = 32'd37243;
			28294: outdata = 32'd37242;
			28295: outdata = 32'd37241;
			28296: outdata = 32'd37240;
			28297: outdata = 32'd37239;
			28298: outdata = 32'd37238;
			28299: outdata = 32'd37237;
			28300: outdata = 32'd37236;
			28301: outdata = 32'd37235;
			28302: outdata = 32'd37234;
			28303: outdata = 32'd37233;
			28304: outdata = 32'd37232;
			28305: outdata = 32'd37231;
			28306: outdata = 32'd37230;
			28307: outdata = 32'd37229;
			28308: outdata = 32'd37228;
			28309: outdata = 32'd37227;
			28310: outdata = 32'd37226;
			28311: outdata = 32'd37225;
			28312: outdata = 32'd37224;
			28313: outdata = 32'd37223;
			28314: outdata = 32'd37222;
			28315: outdata = 32'd37221;
			28316: outdata = 32'd37220;
			28317: outdata = 32'd37219;
			28318: outdata = 32'd37218;
			28319: outdata = 32'd37217;
			28320: outdata = 32'd37216;
			28321: outdata = 32'd37215;
			28322: outdata = 32'd37214;
			28323: outdata = 32'd37213;
			28324: outdata = 32'd37212;
			28325: outdata = 32'd37211;
			28326: outdata = 32'd37210;
			28327: outdata = 32'd37209;
			28328: outdata = 32'd37208;
			28329: outdata = 32'd37207;
			28330: outdata = 32'd37206;
			28331: outdata = 32'd37205;
			28332: outdata = 32'd37204;
			28333: outdata = 32'd37203;
			28334: outdata = 32'd37202;
			28335: outdata = 32'd37201;
			28336: outdata = 32'd37200;
			28337: outdata = 32'd37199;
			28338: outdata = 32'd37198;
			28339: outdata = 32'd37197;
			28340: outdata = 32'd37196;
			28341: outdata = 32'd37195;
			28342: outdata = 32'd37194;
			28343: outdata = 32'd37193;
			28344: outdata = 32'd37192;
			28345: outdata = 32'd37191;
			28346: outdata = 32'd37190;
			28347: outdata = 32'd37189;
			28348: outdata = 32'd37188;
			28349: outdata = 32'd37187;
			28350: outdata = 32'd37186;
			28351: outdata = 32'd37185;
			28352: outdata = 32'd37184;
			28353: outdata = 32'd37183;
			28354: outdata = 32'd37182;
			28355: outdata = 32'd37181;
			28356: outdata = 32'd37180;
			28357: outdata = 32'd37179;
			28358: outdata = 32'd37178;
			28359: outdata = 32'd37177;
			28360: outdata = 32'd37176;
			28361: outdata = 32'd37175;
			28362: outdata = 32'd37174;
			28363: outdata = 32'd37173;
			28364: outdata = 32'd37172;
			28365: outdata = 32'd37171;
			28366: outdata = 32'd37170;
			28367: outdata = 32'd37169;
			28368: outdata = 32'd37168;
			28369: outdata = 32'd37167;
			28370: outdata = 32'd37166;
			28371: outdata = 32'd37165;
			28372: outdata = 32'd37164;
			28373: outdata = 32'd37163;
			28374: outdata = 32'd37162;
			28375: outdata = 32'd37161;
			28376: outdata = 32'd37160;
			28377: outdata = 32'd37159;
			28378: outdata = 32'd37158;
			28379: outdata = 32'd37157;
			28380: outdata = 32'd37156;
			28381: outdata = 32'd37155;
			28382: outdata = 32'd37154;
			28383: outdata = 32'd37153;
			28384: outdata = 32'd37152;
			28385: outdata = 32'd37151;
			28386: outdata = 32'd37150;
			28387: outdata = 32'd37149;
			28388: outdata = 32'd37148;
			28389: outdata = 32'd37147;
			28390: outdata = 32'd37146;
			28391: outdata = 32'd37145;
			28392: outdata = 32'd37144;
			28393: outdata = 32'd37143;
			28394: outdata = 32'd37142;
			28395: outdata = 32'd37141;
			28396: outdata = 32'd37140;
			28397: outdata = 32'd37139;
			28398: outdata = 32'd37138;
			28399: outdata = 32'd37137;
			28400: outdata = 32'd37136;
			28401: outdata = 32'd37135;
			28402: outdata = 32'd37134;
			28403: outdata = 32'd37133;
			28404: outdata = 32'd37132;
			28405: outdata = 32'd37131;
			28406: outdata = 32'd37130;
			28407: outdata = 32'd37129;
			28408: outdata = 32'd37128;
			28409: outdata = 32'd37127;
			28410: outdata = 32'd37126;
			28411: outdata = 32'd37125;
			28412: outdata = 32'd37124;
			28413: outdata = 32'd37123;
			28414: outdata = 32'd37122;
			28415: outdata = 32'd37121;
			28416: outdata = 32'd37120;
			28417: outdata = 32'd37119;
			28418: outdata = 32'd37118;
			28419: outdata = 32'd37117;
			28420: outdata = 32'd37116;
			28421: outdata = 32'd37115;
			28422: outdata = 32'd37114;
			28423: outdata = 32'd37113;
			28424: outdata = 32'd37112;
			28425: outdata = 32'd37111;
			28426: outdata = 32'd37110;
			28427: outdata = 32'd37109;
			28428: outdata = 32'd37108;
			28429: outdata = 32'd37107;
			28430: outdata = 32'd37106;
			28431: outdata = 32'd37105;
			28432: outdata = 32'd37104;
			28433: outdata = 32'd37103;
			28434: outdata = 32'd37102;
			28435: outdata = 32'd37101;
			28436: outdata = 32'd37100;
			28437: outdata = 32'd37099;
			28438: outdata = 32'd37098;
			28439: outdata = 32'd37097;
			28440: outdata = 32'd37096;
			28441: outdata = 32'd37095;
			28442: outdata = 32'd37094;
			28443: outdata = 32'd37093;
			28444: outdata = 32'd37092;
			28445: outdata = 32'd37091;
			28446: outdata = 32'd37090;
			28447: outdata = 32'd37089;
			28448: outdata = 32'd37088;
			28449: outdata = 32'd37087;
			28450: outdata = 32'd37086;
			28451: outdata = 32'd37085;
			28452: outdata = 32'd37084;
			28453: outdata = 32'd37083;
			28454: outdata = 32'd37082;
			28455: outdata = 32'd37081;
			28456: outdata = 32'd37080;
			28457: outdata = 32'd37079;
			28458: outdata = 32'd37078;
			28459: outdata = 32'd37077;
			28460: outdata = 32'd37076;
			28461: outdata = 32'd37075;
			28462: outdata = 32'd37074;
			28463: outdata = 32'd37073;
			28464: outdata = 32'd37072;
			28465: outdata = 32'd37071;
			28466: outdata = 32'd37070;
			28467: outdata = 32'd37069;
			28468: outdata = 32'd37068;
			28469: outdata = 32'd37067;
			28470: outdata = 32'd37066;
			28471: outdata = 32'd37065;
			28472: outdata = 32'd37064;
			28473: outdata = 32'd37063;
			28474: outdata = 32'd37062;
			28475: outdata = 32'd37061;
			28476: outdata = 32'd37060;
			28477: outdata = 32'd37059;
			28478: outdata = 32'd37058;
			28479: outdata = 32'd37057;
			28480: outdata = 32'd37056;
			28481: outdata = 32'd37055;
			28482: outdata = 32'd37054;
			28483: outdata = 32'd37053;
			28484: outdata = 32'd37052;
			28485: outdata = 32'd37051;
			28486: outdata = 32'd37050;
			28487: outdata = 32'd37049;
			28488: outdata = 32'd37048;
			28489: outdata = 32'd37047;
			28490: outdata = 32'd37046;
			28491: outdata = 32'd37045;
			28492: outdata = 32'd37044;
			28493: outdata = 32'd37043;
			28494: outdata = 32'd37042;
			28495: outdata = 32'd37041;
			28496: outdata = 32'd37040;
			28497: outdata = 32'd37039;
			28498: outdata = 32'd37038;
			28499: outdata = 32'd37037;
			28500: outdata = 32'd37036;
			28501: outdata = 32'd37035;
			28502: outdata = 32'd37034;
			28503: outdata = 32'd37033;
			28504: outdata = 32'd37032;
			28505: outdata = 32'd37031;
			28506: outdata = 32'd37030;
			28507: outdata = 32'd37029;
			28508: outdata = 32'd37028;
			28509: outdata = 32'd37027;
			28510: outdata = 32'd37026;
			28511: outdata = 32'd37025;
			28512: outdata = 32'd37024;
			28513: outdata = 32'd37023;
			28514: outdata = 32'd37022;
			28515: outdata = 32'd37021;
			28516: outdata = 32'd37020;
			28517: outdata = 32'd37019;
			28518: outdata = 32'd37018;
			28519: outdata = 32'd37017;
			28520: outdata = 32'd37016;
			28521: outdata = 32'd37015;
			28522: outdata = 32'd37014;
			28523: outdata = 32'd37013;
			28524: outdata = 32'd37012;
			28525: outdata = 32'd37011;
			28526: outdata = 32'd37010;
			28527: outdata = 32'd37009;
			28528: outdata = 32'd37008;
			28529: outdata = 32'd37007;
			28530: outdata = 32'd37006;
			28531: outdata = 32'd37005;
			28532: outdata = 32'd37004;
			28533: outdata = 32'd37003;
			28534: outdata = 32'd37002;
			28535: outdata = 32'd37001;
			28536: outdata = 32'd37000;
			28537: outdata = 32'd36999;
			28538: outdata = 32'd36998;
			28539: outdata = 32'd36997;
			28540: outdata = 32'd36996;
			28541: outdata = 32'd36995;
			28542: outdata = 32'd36994;
			28543: outdata = 32'd36993;
			28544: outdata = 32'd36992;
			28545: outdata = 32'd36991;
			28546: outdata = 32'd36990;
			28547: outdata = 32'd36989;
			28548: outdata = 32'd36988;
			28549: outdata = 32'd36987;
			28550: outdata = 32'd36986;
			28551: outdata = 32'd36985;
			28552: outdata = 32'd36984;
			28553: outdata = 32'd36983;
			28554: outdata = 32'd36982;
			28555: outdata = 32'd36981;
			28556: outdata = 32'd36980;
			28557: outdata = 32'd36979;
			28558: outdata = 32'd36978;
			28559: outdata = 32'd36977;
			28560: outdata = 32'd36976;
			28561: outdata = 32'd36975;
			28562: outdata = 32'd36974;
			28563: outdata = 32'd36973;
			28564: outdata = 32'd36972;
			28565: outdata = 32'd36971;
			28566: outdata = 32'd36970;
			28567: outdata = 32'd36969;
			28568: outdata = 32'd36968;
			28569: outdata = 32'd36967;
			28570: outdata = 32'd36966;
			28571: outdata = 32'd36965;
			28572: outdata = 32'd36964;
			28573: outdata = 32'd36963;
			28574: outdata = 32'd36962;
			28575: outdata = 32'd36961;
			28576: outdata = 32'd36960;
			28577: outdata = 32'd36959;
			28578: outdata = 32'd36958;
			28579: outdata = 32'd36957;
			28580: outdata = 32'd36956;
			28581: outdata = 32'd36955;
			28582: outdata = 32'd36954;
			28583: outdata = 32'd36953;
			28584: outdata = 32'd36952;
			28585: outdata = 32'd36951;
			28586: outdata = 32'd36950;
			28587: outdata = 32'd36949;
			28588: outdata = 32'd36948;
			28589: outdata = 32'd36947;
			28590: outdata = 32'd36946;
			28591: outdata = 32'd36945;
			28592: outdata = 32'd36944;
			28593: outdata = 32'd36943;
			28594: outdata = 32'd36942;
			28595: outdata = 32'd36941;
			28596: outdata = 32'd36940;
			28597: outdata = 32'd36939;
			28598: outdata = 32'd36938;
			28599: outdata = 32'd36937;
			28600: outdata = 32'd36936;
			28601: outdata = 32'd36935;
			28602: outdata = 32'd36934;
			28603: outdata = 32'd36933;
			28604: outdata = 32'd36932;
			28605: outdata = 32'd36931;
			28606: outdata = 32'd36930;
			28607: outdata = 32'd36929;
			28608: outdata = 32'd36928;
			28609: outdata = 32'd36927;
			28610: outdata = 32'd36926;
			28611: outdata = 32'd36925;
			28612: outdata = 32'd36924;
			28613: outdata = 32'd36923;
			28614: outdata = 32'd36922;
			28615: outdata = 32'd36921;
			28616: outdata = 32'd36920;
			28617: outdata = 32'd36919;
			28618: outdata = 32'd36918;
			28619: outdata = 32'd36917;
			28620: outdata = 32'd36916;
			28621: outdata = 32'd36915;
			28622: outdata = 32'd36914;
			28623: outdata = 32'd36913;
			28624: outdata = 32'd36912;
			28625: outdata = 32'd36911;
			28626: outdata = 32'd36910;
			28627: outdata = 32'd36909;
			28628: outdata = 32'd36908;
			28629: outdata = 32'd36907;
			28630: outdata = 32'd36906;
			28631: outdata = 32'd36905;
			28632: outdata = 32'd36904;
			28633: outdata = 32'd36903;
			28634: outdata = 32'd36902;
			28635: outdata = 32'd36901;
			28636: outdata = 32'd36900;
			28637: outdata = 32'd36899;
			28638: outdata = 32'd36898;
			28639: outdata = 32'd36897;
			28640: outdata = 32'd36896;
			28641: outdata = 32'd36895;
			28642: outdata = 32'd36894;
			28643: outdata = 32'd36893;
			28644: outdata = 32'd36892;
			28645: outdata = 32'd36891;
			28646: outdata = 32'd36890;
			28647: outdata = 32'd36889;
			28648: outdata = 32'd36888;
			28649: outdata = 32'd36887;
			28650: outdata = 32'd36886;
			28651: outdata = 32'd36885;
			28652: outdata = 32'd36884;
			28653: outdata = 32'd36883;
			28654: outdata = 32'd36882;
			28655: outdata = 32'd36881;
			28656: outdata = 32'd36880;
			28657: outdata = 32'd36879;
			28658: outdata = 32'd36878;
			28659: outdata = 32'd36877;
			28660: outdata = 32'd36876;
			28661: outdata = 32'd36875;
			28662: outdata = 32'd36874;
			28663: outdata = 32'd36873;
			28664: outdata = 32'd36872;
			28665: outdata = 32'd36871;
			28666: outdata = 32'd36870;
			28667: outdata = 32'd36869;
			28668: outdata = 32'd36868;
			28669: outdata = 32'd36867;
			28670: outdata = 32'd36866;
			28671: outdata = 32'd36865;
			28672: outdata = 32'd36864;
			28673: outdata = 32'd36863;
			28674: outdata = 32'd36862;
			28675: outdata = 32'd36861;
			28676: outdata = 32'd36860;
			28677: outdata = 32'd36859;
			28678: outdata = 32'd36858;
			28679: outdata = 32'd36857;
			28680: outdata = 32'd36856;
			28681: outdata = 32'd36855;
			28682: outdata = 32'd36854;
			28683: outdata = 32'd36853;
			28684: outdata = 32'd36852;
			28685: outdata = 32'd36851;
			28686: outdata = 32'd36850;
			28687: outdata = 32'd36849;
			28688: outdata = 32'd36848;
			28689: outdata = 32'd36847;
			28690: outdata = 32'd36846;
			28691: outdata = 32'd36845;
			28692: outdata = 32'd36844;
			28693: outdata = 32'd36843;
			28694: outdata = 32'd36842;
			28695: outdata = 32'd36841;
			28696: outdata = 32'd36840;
			28697: outdata = 32'd36839;
			28698: outdata = 32'd36838;
			28699: outdata = 32'd36837;
			28700: outdata = 32'd36836;
			28701: outdata = 32'd36835;
			28702: outdata = 32'd36834;
			28703: outdata = 32'd36833;
			28704: outdata = 32'd36832;
			28705: outdata = 32'd36831;
			28706: outdata = 32'd36830;
			28707: outdata = 32'd36829;
			28708: outdata = 32'd36828;
			28709: outdata = 32'd36827;
			28710: outdata = 32'd36826;
			28711: outdata = 32'd36825;
			28712: outdata = 32'd36824;
			28713: outdata = 32'd36823;
			28714: outdata = 32'd36822;
			28715: outdata = 32'd36821;
			28716: outdata = 32'd36820;
			28717: outdata = 32'd36819;
			28718: outdata = 32'd36818;
			28719: outdata = 32'd36817;
			28720: outdata = 32'd36816;
			28721: outdata = 32'd36815;
			28722: outdata = 32'd36814;
			28723: outdata = 32'd36813;
			28724: outdata = 32'd36812;
			28725: outdata = 32'd36811;
			28726: outdata = 32'd36810;
			28727: outdata = 32'd36809;
			28728: outdata = 32'd36808;
			28729: outdata = 32'd36807;
			28730: outdata = 32'd36806;
			28731: outdata = 32'd36805;
			28732: outdata = 32'd36804;
			28733: outdata = 32'd36803;
			28734: outdata = 32'd36802;
			28735: outdata = 32'd36801;
			28736: outdata = 32'd36800;
			28737: outdata = 32'd36799;
			28738: outdata = 32'd36798;
			28739: outdata = 32'd36797;
			28740: outdata = 32'd36796;
			28741: outdata = 32'd36795;
			28742: outdata = 32'd36794;
			28743: outdata = 32'd36793;
			28744: outdata = 32'd36792;
			28745: outdata = 32'd36791;
			28746: outdata = 32'd36790;
			28747: outdata = 32'd36789;
			28748: outdata = 32'd36788;
			28749: outdata = 32'd36787;
			28750: outdata = 32'd36786;
			28751: outdata = 32'd36785;
			28752: outdata = 32'd36784;
			28753: outdata = 32'd36783;
			28754: outdata = 32'd36782;
			28755: outdata = 32'd36781;
			28756: outdata = 32'd36780;
			28757: outdata = 32'd36779;
			28758: outdata = 32'd36778;
			28759: outdata = 32'd36777;
			28760: outdata = 32'd36776;
			28761: outdata = 32'd36775;
			28762: outdata = 32'd36774;
			28763: outdata = 32'd36773;
			28764: outdata = 32'd36772;
			28765: outdata = 32'd36771;
			28766: outdata = 32'd36770;
			28767: outdata = 32'd36769;
			28768: outdata = 32'd36768;
			28769: outdata = 32'd36767;
			28770: outdata = 32'd36766;
			28771: outdata = 32'd36765;
			28772: outdata = 32'd36764;
			28773: outdata = 32'd36763;
			28774: outdata = 32'd36762;
			28775: outdata = 32'd36761;
			28776: outdata = 32'd36760;
			28777: outdata = 32'd36759;
			28778: outdata = 32'd36758;
			28779: outdata = 32'd36757;
			28780: outdata = 32'd36756;
			28781: outdata = 32'd36755;
			28782: outdata = 32'd36754;
			28783: outdata = 32'd36753;
			28784: outdata = 32'd36752;
			28785: outdata = 32'd36751;
			28786: outdata = 32'd36750;
			28787: outdata = 32'd36749;
			28788: outdata = 32'd36748;
			28789: outdata = 32'd36747;
			28790: outdata = 32'd36746;
			28791: outdata = 32'd36745;
			28792: outdata = 32'd36744;
			28793: outdata = 32'd36743;
			28794: outdata = 32'd36742;
			28795: outdata = 32'd36741;
			28796: outdata = 32'd36740;
			28797: outdata = 32'd36739;
			28798: outdata = 32'd36738;
			28799: outdata = 32'd36737;
			28800: outdata = 32'd36736;
			28801: outdata = 32'd36735;
			28802: outdata = 32'd36734;
			28803: outdata = 32'd36733;
			28804: outdata = 32'd36732;
			28805: outdata = 32'd36731;
			28806: outdata = 32'd36730;
			28807: outdata = 32'd36729;
			28808: outdata = 32'd36728;
			28809: outdata = 32'd36727;
			28810: outdata = 32'd36726;
			28811: outdata = 32'd36725;
			28812: outdata = 32'd36724;
			28813: outdata = 32'd36723;
			28814: outdata = 32'd36722;
			28815: outdata = 32'd36721;
			28816: outdata = 32'd36720;
			28817: outdata = 32'd36719;
			28818: outdata = 32'd36718;
			28819: outdata = 32'd36717;
			28820: outdata = 32'd36716;
			28821: outdata = 32'd36715;
			28822: outdata = 32'd36714;
			28823: outdata = 32'd36713;
			28824: outdata = 32'd36712;
			28825: outdata = 32'd36711;
			28826: outdata = 32'd36710;
			28827: outdata = 32'd36709;
			28828: outdata = 32'd36708;
			28829: outdata = 32'd36707;
			28830: outdata = 32'd36706;
			28831: outdata = 32'd36705;
			28832: outdata = 32'd36704;
			28833: outdata = 32'd36703;
			28834: outdata = 32'd36702;
			28835: outdata = 32'd36701;
			28836: outdata = 32'd36700;
			28837: outdata = 32'd36699;
			28838: outdata = 32'd36698;
			28839: outdata = 32'd36697;
			28840: outdata = 32'd36696;
			28841: outdata = 32'd36695;
			28842: outdata = 32'd36694;
			28843: outdata = 32'd36693;
			28844: outdata = 32'd36692;
			28845: outdata = 32'd36691;
			28846: outdata = 32'd36690;
			28847: outdata = 32'd36689;
			28848: outdata = 32'd36688;
			28849: outdata = 32'd36687;
			28850: outdata = 32'd36686;
			28851: outdata = 32'd36685;
			28852: outdata = 32'd36684;
			28853: outdata = 32'd36683;
			28854: outdata = 32'd36682;
			28855: outdata = 32'd36681;
			28856: outdata = 32'd36680;
			28857: outdata = 32'd36679;
			28858: outdata = 32'd36678;
			28859: outdata = 32'd36677;
			28860: outdata = 32'd36676;
			28861: outdata = 32'd36675;
			28862: outdata = 32'd36674;
			28863: outdata = 32'd36673;
			28864: outdata = 32'd36672;
			28865: outdata = 32'd36671;
			28866: outdata = 32'd36670;
			28867: outdata = 32'd36669;
			28868: outdata = 32'd36668;
			28869: outdata = 32'd36667;
			28870: outdata = 32'd36666;
			28871: outdata = 32'd36665;
			28872: outdata = 32'd36664;
			28873: outdata = 32'd36663;
			28874: outdata = 32'd36662;
			28875: outdata = 32'd36661;
			28876: outdata = 32'd36660;
			28877: outdata = 32'd36659;
			28878: outdata = 32'd36658;
			28879: outdata = 32'd36657;
			28880: outdata = 32'd36656;
			28881: outdata = 32'd36655;
			28882: outdata = 32'd36654;
			28883: outdata = 32'd36653;
			28884: outdata = 32'd36652;
			28885: outdata = 32'd36651;
			28886: outdata = 32'd36650;
			28887: outdata = 32'd36649;
			28888: outdata = 32'd36648;
			28889: outdata = 32'd36647;
			28890: outdata = 32'd36646;
			28891: outdata = 32'd36645;
			28892: outdata = 32'd36644;
			28893: outdata = 32'd36643;
			28894: outdata = 32'd36642;
			28895: outdata = 32'd36641;
			28896: outdata = 32'd36640;
			28897: outdata = 32'd36639;
			28898: outdata = 32'd36638;
			28899: outdata = 32'd36637;
			28900: outdata = 32'd36636;
			28901: outdata = 32'd36635;
			28902: outdata = 32'd36634;
			28903: outdata = 32'd36633;
			28904: outdata = 32'd36632;
			28905: outdata = 32'd36631;
			28906: outdata = 32'd36630;
			28907: outdata = 32'd36629;
			28908: outdata = 32'd36628;
			28909: outdata = 32'd36627;
			28910: outdata = 32'd36626;
			28911: outdata = 32'd36625;
			28912: outdata = 32'd36624;
			28913: outdata = 32'd36623;
			28914: outdata = 32'd36622;
			28915: outdata = 32'd36621;
			28916: outdata = 32'd36620;
			28917: outdata = 32'd36619;
			28918: outdata = 32'd36618;
			28919: outdata = 32'd36617;
			28920: outdata = 32'd36616;
			28921: outdata = 32'd36615;
			28922: outdata = 32'd36614;
			28923: outdata = 32'd36613;
			28924: outdata = 32'd36612;
			28925: outdata = 32'd36611;
			28926: outdata = 32'd36610;
			28927: outdata = 32'd36609;
			28928: outdata = 32'd36608;
			28929: outdata = 32'd36607;
			28930: outdata = 32'd36606;
			28931: outdata = 32'd36605;
			28932: outdata = 32'd36604;
			28933: outdata = 32'd36603;
			28934: outdata = 32'd36602;
			28935: outdata = 32'd36601;
			28936: outdata = 32'd36600;
			28937: outdata = 32'd36599;
			28938: outdata = 32'd36598;
			28939: outdata = 32'd36597;
			28940: outdata = 32'd36596;
			28941: outdata = 32'd36595;
			28942: outdata = 32'd36594;
			28943: outdata = 32'd36593;
			28944: outdata = 32'd36592;
			28945: outdata = 32'd36591;
			28946: outdata = 32'd36590;
			28947: outdata = 32'd36589;
			28948: outdata = 32'd36588;
			28949: outdata = 32'd36587;
			28950: outdata = 32'd36586;
			28951: outdata = 32'd36585;
			28952: outdata = 32'd36584;
			28953: outdata = 32'd36583;
			28954: outdata = 32'd36582;
			28955: outdata = 32'd36581;
			28956: outdata = 32'd36580;
			28957: outdata = 32'd36579;
			28958: outdata = 32'd36578;
			28959: outdata = 32'd36577;
			28960: outdata = 32'd36576;
			28961: outdata = 32'd36575;
			28962: outdata = 32'd36574;
			28963: outdata = 32'd36573;
			28964: outdata = 32'd36572;
			28965: outdata = 32'd36571;
			28966: outdata = 32'd36570;
			28967: outdata = 32'd36569;
			28968: outdata = 32'd36568;
			28969: outdata = 32'd36567;
			28970: outdata = 32'd36566;
			28971: outdata = 32'd36565;
			28972: outdata = 32'd36564;
			28973: outdata = 32'd36563;
			28974: outdata = 32'd36562;
			28975: outdata = 32'd36561;
			28976: outdata = 32'd36560;
			28977: outdata = 32'd36559;
			28978: outdata = 32'd36558;
			28979: outdata = 32'd36557;
			28980: outdata = 32'd36556;
			28981: outdata = 32'd36555;
			28982: outdata = 32'd36554;
			28983: outdata = 32'd36553;
			28984: outdata = 32'd36552;
			28985: outdata = 32'd36551;
			28986: outdata = 32'd36550;
			28987: outdata = 32'd36549;
			28988: outdata = 32'd36548;
			28989: outdata = 32'd36547;
			28990: outdata = 32'd36546;
			28991: outdata = 32'd36545;
			28992: outdata = 32'd36544;
			28993: outdata = 32'd36543;
			28994: outdata = 32'd36542;
			28995: outdata = 32'd36541;
			28996: outdata = 32'd36540;
			28997: outdata = 32'd36539;
			28998: outdata = 32'd36538;
			28999: outdata = 32'd36537;
			29000: outdata = 32'd36536;
			29001: outdata = 32'd36535;
			29002: outdata = 32'd36534;
			29003: outdata = 32'd36533;
			29004: outdata = 32'd36532;
			29005: outdata = 32'd36531;
			29006: outdata = 32'd36530;
			29007: outdata = 32'd36529;
			29008: outdata = 32'd36528;
			29009: outdata = 32'd36527;
			29010: outdata = 32'd36526;
			29011: outdata = 32'd36525;
			29012: outdata = 32'd36524;
			29013: outdata = 32'd36523;
			29014: outdata = 32'd36522;
			29015: outdata = 32'd36521;
			29016: outdata = 32'd36520;
			29017: outdata = 32'd36519;
			29018: outdata = 32'd36518;
			29019: outdata = 32'd36517;
			29020: outdata = 32'd36516;
			29021: outdata = 32'd36515;
			29022: outdata = 32'd36514;
			29023: outdata = 32'd36513;
			29024: outdata = 32'd36512;
			29025: outdata = 32'd36511;
			29026: outdata = 32'd36510;
			29027: outdata = 32'd36509;
			29028: outdata = 32'd36508;
			29029: outdata = 32'd36507;
			29030: outdata = 32'd36506;
			29031: outdata = 32'd36505;
			29032: outdata = 32'd36504;
			29033: outdata = 32'd36503;
			29034: outdata = 32'd36502;
			29035: outdata = 32'd36501;
			29036: outdata = 32'd36500;
			29037: outdata = 32'd36499;
			29038: outdata = 32'd36498;
			29039: outdata = 32'd36497;
			29040: outdata = 32'd36496;
			29041: outdata = 32'd36495;
			29042: outdata = 32'd36494;
			29043: outdata = 32'd36493;
			29044: outdata = 32'd36492;
			29045: outdata = 32'd36491;
			29046: outdata = 32'd36490;
			29047: outdata = 32'd36489;
			29048: outdata = 32'd36488;
			29049: outdata = 32'd36487;
			29050: outdata = 32'd36486;
			29051: outdata = 32'd36485;
			29052: outdata = 32'd36484;
			29053: outdata = 32'd36483;
			29054: outdata = 32'd36482;
			29055: outdata = 32'd36481;
			29056: outdata = 32'd36480;
			29057: outdata = 32'd36479;
			29058: outdata = 32'd36478;
			29059: outdata = 32'd36477;
			29060: outdata = 32'd36476;
			29061: outdata = 32'd36475;
			29062: outdata = 32'd36474;
			29063: outdata = 32'd36473;
			29064: outdata = 32'd36472;
			29065: outdata = 32'd36471;
			29066: outdata = 32'd36470;
			29067: outdata = 32'd36469;
			29068: outdata = 32'd36468;
			29069: outdata = 32'd36467;
			29070: outdata = 32'd36466;
			29071: outdata = 32'd36465;
			29072: outdata = 32'd36464;
			29073: outdata = 32'd36463;
			29074: outdata = 32'd36462;
			29075: outdata = 32'd36461;
			29076: outdata = 32'd36460;
			29077: outdata = 32'd36459;
			29078: outdata = 32'd36458;
			29079: outdata = 32'd36457;
			29080: outdata = 32'd36456;
			29081: outdata = 32'd36455;
			29082: outdata = 32'd36454;
			29083: outdata = 32'd36453;
			29084: outdata = 32'd36452;
			29085: outdata = 32'd36451;
			29086: outdata = 32'd36450;
			29087: outdata = 32'd36449;
			29088: outdata = 32'd36448;
			29089: outdata = 32'd36447;
			29090: outdata = 32'd36446;
			29091: outdata = 32'd36445;
			29092: outdata = 32'd36444;
			29093: outdata = 32'd36443;
			29094: outdata = 32'd36442;
			29095: outdata = 32'd36441;
			29096: outdata = 32'd36440;
			29097: outdata = 32'd36439;
			29098: outdata = 32'd36438;
			29099: outdata = 32'd36437;
			29100: outdata = 32'd36436;
			29101: outdata = 32'd36435;
			29102: outdata = 32'd36434;
			29103: outdata = 32'd36433;
			29104: outdata = 32'd36432;
			29105: outdata = 32'd36431;
			29106: outdata = 32'd36430;
			29107: outdata = 32'd36429;
			29108: outdata = 32'd36428;
			29109: outdata = 32'd36427;
			29110: outdata = 32'd36426;
			29111: outdata = 32'd36425;
			29112: outdata = 32'd36424;
			29113: outdata = 32'd36423;
			29114: outdata = 32'd36422;
			29115: outdata = 32'd36421;
			29116: outdata = 32'd36420;
			29117: outdata = 32'd36419;
			29118: outdata = 32'd36418;
			29119: outdata = 32'd36417;
			29120: outdata = 32'd36416;
			29121: outdata = 32'd36415;
			29122: outdata = 32'd36414;
			29123: outdata = 32'd36413;
			29124: outdata = 32'd36412;
			29125: outdata = 32'd36411;
			29126: outdata = 32'd36410;
			29127: outdata = 32'd36409;
			29128: outdata = 32'd36408;
			29129: outdata = 32'd36407;
			29130: outdata = 32'd36406;
			29131: outdata = 32'd36405;
			29132: outdata = 32'd36404;
			29133: outdata = 32'd36403;
			29134: outdata = 32'd36402;
			29135: outdata = 32'd36401;
			29136: outdata = 32'd36400;
			29137: outdata = 32'd36399;
			29138: outdata = 32'd36398;
			29139: outdata = 32'd36397;
			29140: outdata = 32'd36396;
			29141: outdata = 32'd36395;
			29142: outdata = 32'd36394;
			29143: outdata = 32'd36393;
			29144: outdata = 32'd36392;
			29145: outdata = 32'd36391;
			29146: outdata = 32'd36390;
			29147: outdata = 32'd36389;
			29148: outdata = 32'd36388;
			29149: outdata = 32'd36387;
			29150: outdata = 32'd36386;
			29151: outdata = 32'd36385;
			29152: outdata = 32'd36384;
			29153: outdata = 32'd36383;
			29154: outdata = 32'd36382;
			29155: outdata = 32'd36381;
			29156: outdata = 32'd36380;
			29157: outdata = 32'd36379;
			29158: outdata = 32'd36378;
			29159: outdata = 32'd36377;
			29160: outdata = 32'd36376;
			29161: outdata = 32'd36375;
			29162: outdata = 32'd36374;
			29163: outdata = 32'd36373;
			29164: outdata = 32'd36372;
			29165: outdata = 32'd36371;
			29166: outdata = 32'd36370;
			29167: outdata = 32'd36369;
			29168: outdata = 32'd36368;
			29169: outdata = 32'd36367;
			29170: outdata = 32'd36366;
			29171: outdata = 32'd36365;
			29172: outdata = 32'd36364;
			29173: outdata = 32'd36363;
			29174: outdata = 32'd36362;
			29175: outdata = 32'd36361;
			29176: outdata = 32'd36360;
			29177: outdata = 32'd36359;
			29178: outdata = 32'd36358;
			29179: outdata = 32'd36357;
			29180: outdata = 32'd36356;
			29181: outdata = 32'd36355;
			29182: outdata = 32'd36354;
			29183: outdata = 32'd36353;
			29184: outdata = 32'd36352;
			29185: outdata = 32'd36351;
			29186: outdata = 32'd36350;
			29187: outdata = 32'd36349;
			29188: outdata = 32'd36348;
			29189: outdata = 32'd36347;
			29190: outdata = 32'd36346;
			29191: outdata = 32'd36345;
			29192: outdata = 32'd36344;
			29193: outdata = 32'd36343;
			29194: outdata = 32'd36342;
			29195: outdata = 32'd36341;
			29196: outdata = 32'd36340;
			29197: outdata = 32'd36339;
			29198: outdata = 32'd36338;
			29199: outdata = 32'd36337;
			29200: outdata = 32'd36336;
			29201: outdata = 32'd36335;
			29202: outdata = 32'd36334;
			29203: outdata = 32'd36333;
			29204: outdata = 32'd36332;
			29205: outdata = 32'd36331;
			29206: outdata = 32'd36330;
			29207: outdata = 32'd36329;
			29208: outdata = 32'd36328;
			29209: outdata = 32'd36327;
			29210: outdata = 32'd36326;
			29211: outdata = 32'd36325;
			29212: outdata = 32'd36324;
			29213: outdata = 32'd36323;
			29214: outdata = 32'd36322;
			29215: outdata = 32'd36321;
			29216: outdata = 32'd36320;
			29217: outdata = 32'd36319;
			29218: outdata = 32'd36318;
			29219: outdata = 32'd36317;
			29220: outdata = 32'd36316;
			29221: outdata = 32'd36315;
			29222: outdata = 32'd36314;
			29223: outdata = 32'd36313;
			29224: outdata = 32'd36312;
			29225: outdata = 32'd36311;
			29226: outdata = 32'd36310;
			29227: outdata = 32'd36309;
			29228: outdata = 32'd36308;
			29229: outdata = 32'd36307;
			29230: outdata = 32'd36306;
			29231: outdata = 32'd36305;
			29232: outdata = 32'd36304;
			29233: outdata = 32'd36303;
			29234: outdata = 32'd36302;
			29235: outdata = 32'd36301;
			29236: outdata = 32'd36300;
			29237: outdata = 32'd36299;
			29238: outdata = 32'd36298;
			29239: outdata = 32'd36297;
			29240: outdata = 32'd36296;
			29241: outdata = 32'd36295;
			29242: outdata = 32'd36294;
			29243: outdata = 32'd36293;
			29244: outdata = 32'd36292;
			29245: outdata = 32'd36291;
			29246: outdata = 32'd36290;
			29247: outdata = 32'd36289;
			29248: outdata = 32'd36288;
			29249: outdata = 32'd36287;
			29250: outdata = 32'd36286;
			29251: outdata = 32'd36285;
			29252: outdata = 32'd36284;
			29253: outdata = 32'd36283;
			29254: outdata = 32'd36282;
			29255: outdata = 32'd36281;
			29256: outdata = 32'd36280;
			29257: outdata = 32'd36279;
			29258: outdata = 32'd36278;
			29259: outdata = 32'd36277;
			29260: outdata = 32'd36276;
			29261: outdata = 32'd36275;
			29262: outdata = 32'd36274;
			29263: outdata = 32'd36273;
			29264: outdata = 32'd36272;
			29265: outdata = 32'd36271;
			29266: outdata = 32'd36270;
			29267: outdata = 32'd36269;
			29268: outdata = 32'd36268;
			29269: outdata = 32'd36267;
			29270: outdata = 32'd36266;
			29271: outdata = 32'd36265;
			29272: outdata = 32'd36264;
			29273: outdata = 32'd36263;
			29274: outdata = 32'd36262;
			29275: outdata = 32'd36261;
			29276: outdata = 32'd36260;
			29277: outdata = 32'd36259;
			29278: outdata = 32'd36258;
			29279: outdata = 32'd36257;
			29280: outdata = 32'd36256;
			29281: outdata = 32'd36255;
			29282: outdata = 32'd36254;
			29283: outdata = 32'd36253;
			29284: outdata = 32'd36252;
			29285: outdata = 32'd36251;
			29286: outdata = 32'd36250;
			29287: outdata = 32'd36249;
			29288: outdata = 32'd36248;
			29289: outdata = 32'd36247;
			29290: outdata = 32'd36246;
			29291: outdata = 32'd36245;
			29292: outdata = 32'd36244;
			29293: outdata = 32'd36243;
			29294: outdata = 32'd36242;
			29295: outdata = 32'd36241;
			29296: outdata = 32'd36240;
			29297: outdata = 32'd36239;
			29298: outdata = 32'd36238;
			29299: outdata = 32'd36237;
			29300: outdata = 32'd36236;
			29301: outdata = 32'd36235;
			29302: outdata = 32'd36234;
			29303: outdata = 32'd36233;
			29304: outdata = 32'd36232;
			29305: outdata = 32'd36231;
			29306: outdata = 32'd36230;
			29307: outdata = 32'd36229;
			29308: outdata = 32'd36228;
			29309: outdata = 32'd36227;
			29310: outdata = 32'd36226;
			29311: outdata = 32'd36225;
			29312: outdata = 32'd36224;
			29313: outdata = 32'd36223;
			29314: outdata = 32'd36222;
			29315: outdata = 32'd36221;
			29316: outdata = 32'd36220;
			29317: outdata = 32'd36219;
			29318: outdata = 32'd36218;
			29319: outdata = 32'd36217;
			29320: outdata = 32'd36216;
			29321: outdata = 32'd36215;
			29322: outdata = 32'd36214;
			29323: outdata = 32'd36213;
			29324: outdata = 32'd36212;
			29325: outdata = 32'd36211;
			29326: outdata = 32'd36210;
			29327: outdata = 32'd36209;
			29328: outdata = 32'd36208;
			29329: outdata = 32'd36207;
			29330: outdata = 32'd36206;
			29331: outdata = 32'd36205;
			29332: outdata = 32'd36204;
			29333: outdata = 32'd36203;
			29334: outdata = 32'd36202;
			29335: outdata = 32'd36201;
			29336: outdata = 32'd36200;
			29337: outdata = 32'd36199;
			29338: outdata = 32'd36198;
			29339: outdata = 32'd36197;
			29340: outdata = 32'd36196;
			29341: outdata = 32'd36195;
			29342: outdata = 32'd36194;
			29343: outdata = 32'd36193;
			29344: outdata = 32'd36192;
			29345: outdata = 32'd36191;
			29346: outdata = 32'd36190;
			29347: outdata = 32'd36189;
			29348: outdata = 32'd36188;
			29349: outdata = 32'd36187;
			29350: outdata = 32'd36186;
			29351: outdata = 32'd36185;
			29352: outdata = 32'd36184;
			29353: outdata = 32'd36183;
			29354: outdata = 32'd36182;
			29355: outdata = 32'd36181;
			29356: outdata = 32'd36180;
			29357: outdata = 32'd36179;
			29358: outdata = 32'd36178;
			29359: outdata = 32'd36177;
			29360: outdata = 32'd36176;
			29361: outdata = 32'd36175;
			29362: outdata = 32'd36174;
			29363: outdata = 32'd36173;
			29364: outdata = 32'd36172;
			29365: outdata = 32'd36171;
			29366: outdata = 32'd36170;
			29367: outdata = 32'd36169;
			29368: outdata = 32'd36168;
			29369: outdata = 32'd36167;
			29370: outdata = 32'd36166;
			29371: outdata = 32'd36165;
			29372: outdata = 32'd36164;
			29373: outdata = 32'd36163;
			29374: outdata = 32'd36162;
			29375: outdata = 32'd36161;
			29376: outdata = 32'd36160;
			29377: outdata = 32'd36159;
			29378: outdata = 32'd36158;
			29379: outdata = 32'd36157;
			29380: outdata = 32'd36156;
			29381: outdata = 32'd36155;
			29382: outdata = 32'd36154;
			29383: outdata = 32'd36153;
			29384: outdata = 32'd36152;
			29385: outdata = 32'd36151;
			29386: outdata = 32'd36150;
			29387: outdata = 32'd36149;
			29388: outdata = 32'd36148;
			29389: outdata = 32'd36147;
			29390: outdata = 32'd36146;
			29391: outdata = 32'd36145;
			29392: outdata = 32'd36144;
			29393: outdata = 32'd36143;
			29394: outdata = 32'd36142;
			29395: outdata = 32'd36141;
			29396: outdata = 32'd36140;
			29397: outdata = 32'd36139;
			29398: outdata = 32'd36138;
			29399: outdata = 32'd36137;
			29400: outdata = 32'd36136;
			29401: outdata = 32'd36135;
			29402: outdata = 32'd36134;
			29403: outdata = 32'd36133;
			29404: outdata = 32'd36132;
			29405: outdata = 32'd36131;
			29406: outdata = 32'd36130;
			29407: outdata = 32'd36129;
			29408: outdata = 32'd36128;
			29409: outdata = 32'd36127;
			29410: outdata = 32'd36126;
			29411: outdata = 32'd36125;
			29412: outdata = 32'd36124;
			29413: outdata = 32'd36123;
			29414: outdata = 32'd36122;
			29415: outdata = 32'd36121;
			29416: outdata = 32'd36120;
			29417: outdata = 32'd36119;
			29418: outdata = 32'd36118;
			29419: outdata = 32'd36117;
			29420: outdata = 32'd36116;
			29421: outdata = 32'd36115;
			29422: outdata = 32'd36114;
			29423: outdata = 32'd36113;
			29424: outdata = 32'd36112;
			29425: outdata = 32'd36111;
			29426: outdata = 32'd36110;
			29427: outdata = 32'd36109;
			29428: outdata = 32'd36108;
			29429: outdata = 32'd36107;
			29430: outdata = 32'd36106;
			29431: outdata = 32'd36105;
			29432: outdata = 32'd36104;
			29433: outdata = 32'd36103;
			29434: outdata = 32'd36102;
			29435: outdata = 32'd36101;
			29436: outdata = 32'd36100;
			29437: outdata = 32'd36099;
			29438: outdata = 32'd36098;
			29439: outdata = 32'd36097;
			29440: outdata = 32'd36096;
			29441: outdata = 32'd36095;
			29442: outdata = 32'd36094;
			29443: outdata = 32'd36093;
			29444: outdata = 32'd36092;
			29445: outdata = 32'd36091;
			29446: outdata = 32'd36090;
			29447: outdata = 32'd36089;
			29448: outdata = 32'd36088;
			29449: outdata = 32'd36087;
			29450: outdata = 32'd36086;
			29451: outdata = 32'd36085;
			29452: outdata = 32'd36084;
			29453: outdata = 32'd36083;
			29454: outdata = 32'd36082;
			29455: outdata = 32'd36081;
			29456: outdata = 32'd36080;
			29457: outdata = 32'd36079;
			29458: outdata = 32'd36078;
			29459: outdata = 32'd36077;
			29460: outdata = 32'd36076;
			29461: outdata = 32'd36075;
			29462: outdata = 32'd36074;
			29463: outdata = 32'd36073;
			29464: outdata = 32'd36072;
			29465: outdata = 32'd36071;
			29466: outdata = 32'd36070;
			29467: outdata = 32'd36069;
			29468: outdata = 32'd36068;
			29469: outdata = 32'd36067;
			29470: outdata = 32'd36066;
			29471: outdata = 32'd36065;
			29472: outdata = 32'd36064;
			29473: outdata = 32'd36063;
			29474: outdata = 32'd36062;
			29475: outdata = 32'd36061;
			29476: outdata = 32'd36060;
			29477: outdata = 32'd36059;
			29478: outdata = 32'd36058;
			29479: outdata = 32'd36057;
			29480: outdata = 32'd36056;
			29481: outdata = 32'd36055;
			29482: outdata = 32'd36054;
			29483: outdata = 32'd36053;
			29484: outdata = 32'd36052;
			29485: outdata = 32'd36051;
			29486: outdata = 32'd36050;
			29487: outdata = 32'd36049;
			29488: outdata = 32'd36048;
			29489: outdata = 32'd36047;
			29490: outdata = 32'd36046;
			29491: outdata = 32'd36045;
			29492: outdata = 32'd36044;
			29493: outdata = 32'd36043;
			29494: outdata = 32'd36042;
			29495: outdata = 32'd36041;
			29496: outdata = 32'd36040;
			29497: outdata = 32'd36039;
			29498: outdata = 32'd36038;
			29499: outdata = 32'd36037;
			29500: outdata = 32'd36036;
			29501: outdata = 32'd36035;
			29502: outdata = 32'd36034;
			29503: outdata = 32'd36033;
			29504: outdata = 32'd36032;
			29505: outdata = 32'd36031;
			29506: outdata = 32'd36030;
			29507: outdata = 32'd36029;
			29508: outdata = 32'd36028;
			29509: outdata = 32'd36027;
			29510: outdata = 32'd36026;
			29511: outdata = 32'd36025;
			29512: outdata = 32'd36024;
			29513: outdata = 32'd36023;
			29514: outdata = 32'd36022;
			29515: outdata = 32'd36021;
			29516: outdata = 32'd36020;
			29517: outdata = 32'd36019;
			29518: outdata = 32'd36018;
			29519: outdata = 32'd36017;
			29520: outdata = 32'd36016;
			29521: outdata = 32'd36015;
			29522: outdata = 32'd36014;
			29523: outdata = 32'd36013;
			29524: outdata = 32'd36012;
			29525: outdata = 32'd36011;
			29526: outdata = 32'd36010;
			29527: outdata = 32'd36009;
			29528: outdata = 32'd36008;
			29529: outdata = 32'd36007;
			29530: outdata = 32'd36006;
			29531: outdata = 32'd36005;
			29532: outdata = 32'd36004;
			29533: outdata = 32'd36003;
			29534: outdata = 32'd36002;
			29535: outdata = 32'd36001;
			29536: outdata = 32'd36000;
			29537: outdata = 32'd35999;
			29538: outdata = 32'd35998;
			29539: outdata = 32'd35997;
			29540: outdata = 32'd35996;
			29541: outdata = 32'd35995;
			29542: outdata = 32'd35994;
			29543: outdata = 32'd35993;
			29544: outdata = 32'd35992;
			29545: outdata = 32'd35991;
			29546: outdata = 32'd35990;
			29547: outdata = 32'd35989;
			29548: outdata = 32'd35988;
			29549: outdata = 32'd35987;
			29550: outdata = 32'd35986;
			29551: outdata = 32'd35985;
			29552: outdata = 32'd35984;
			29553: outdata = 32'd35983;
			29554: outdata = 32'd35982;
			29555: outdata = 32'd35981;
			29556: outdata = 32'd35980;
			29557: outdata = 32'd35979;
			29558: outdata = 32'd35978;
			29559: outdata = 32'd35977;
			29560: outdata = 32'd35976;
			29561: outdata = 32'd35975;
			29562: outdata = 32'd35974;
			29563: outdata = 32'd35973;
			29564: outdata = 32'd35972;
			29565: outdata = 32'd35971;
			29566: outdata = 32'd35970;
			29567: outdata = 32'd35969;
			29568: outdata = 32'd35968;
			29569: outdata = 32'd35967;
			29570: outdata = 32'd35966;
			29571: outdata = 32'd35965;
			29572: outdata = 32'd35964;
			29573: outdata = 32'd35963;
			29574: outdata = 32'd35962;
			29575: outdata = 32'd35961;
			29576: outdata = 32'd35960;
			29577: outdata = 32'd35959;
			29578: outdata = 32'd35958;
			29579: outdata = 32'd35957;
			29580: outdata = 32'd35956;
			29581: outdata = 32'd35955;
			29582: outdata = 32'd35954;
			29583: outdata = 32'd35953;
			29584: outdata = 32'd35952;
			29585: outdata = 32'd35951;
			29586: outdata = 32'd35950;
			29587: outdata = 32'd35949;
			29588: outdata = 32'd35948;
			29589: outdata = 32'd35947;
			29590: outdata = 32'd35946;
			29591: outdata = 32'd35945;
			29592: outdata = 32'd35944;
			29593: outdata = 32'd35943;
			29594: outdata = 32'd35942;
			29595: outdata = 32'd35941;
			29596: outdata = 32'd35940;
			29597: outdata = 32'd35939;
			29598: outdata = 32'd35938;
			29599: outdata = 32'd35937;
			29600: outdata = 32'd35936;
			29601: outdata = 32'd35935;
			29602: outdata = 32'd35934;
			29603: outdata = 32'd35933;
			29604: outdata = 32'd35932;
			29605: outdata = 32'd35931;
			29606: outdata = 32'd35930;
			29607: outdata = 32'd35929;
			29608: outdata = 32'd35928;
			29609: outdata = 32'd35927;
			29610: outdata = 32'd35926;
			29611: outdata = 32'd35925;
			29612: outdata = 32'd35924;
			29613: outdata = 32'd35923;
			29614: outdata = 32'd35922;
			29615: outdata = 32'd35921;
			29616: outdata = 32'd35920;
			29617: outdata = 32'd35919;
			29618: outdata = 32'd35918;
			29619: outdata = 32'd35917;
			29620: outdata = 32'd35916;
			29621: outdata = 32'd35915;
			29622: outdata = 32'd35914;
			29623: outdata = 32'd35913;
			29624: outdata = 32'd35912;
			29625: outdata = 32'd35911;
			29626: outdata = 32'd35910;
			29627: outdata = 32'd35909;
			29628: outdata = 32'd35908;
			29629: outdata = 32'd35907;
			29630: outdata = 32'd35906;
			29631: outdata = 32'd35905;
			29632: outdata = 32'd35904;
			29633: outdata = 32'd35903;
			29634: outdata = 32'd35902;
			29635: outdata = 32'd35901;
			29636: outdata = 32'd35900;
			29637: outdata = 32'd35899;
			29638: outdata = 32'd35898;
			29639: outdata = 32'd35897;
			29640: outdata = 32'd35896;
			29641: outdata = 32'd35895;
			29642: outdata = 32'd35894;
			29643: outdata = 32'd35893;
			29644: outdata = 32'd35892;
			29645: outdata = 32'd35891;
			29646: outdata = 32'd35890;
			29647: outdata = 32'd35889;
			29648: outdata = 32'd35888;
			29649: outdata = 32'd35887;
			29650: outdata = 32'd35886;
			29651: outdata = 32'd35885;
			29652: outdata = 32'd35884;
			29653: outdata = 32'd35883;
			29654: outdata = 32'd35882;
			29655: outdata = 32'd35881;
			29656: outdata = 32'd35880;
			29657: outdata = 32'd35879;
			29658: outdata = 32'd35878;
			29659: outdata = 32'd35877;
			29660: outdata = 32'd35876;
			29661: outdata = 32'd35875;
			29662: outdata = 32'd35874;
			29663: outdata = 32'd35873;
			29664: outdata = 32'd35872;
			29665: outdata = 32'd35871;
			29666: outdata = 32'd35870;
			29667: outdata = 32'd35869;
			29668: outdata = 32'd35868;
			29669: outdata = 32'd35867;
			29670: outdata = 32'd35866;
			29671: outdata = 32'd35865;
			29672: outdata = 32'd35864;
			29673: outdata = 32'd35863;
			29674: outdata = 32'd35862;
			29675: outdata = 32'd35861;
			29676: outdata = 32'd35860;
			29677: outdata = 32'd35859;
			29678: outdata = 32'd35858;
			29679: outdata = 32'd35857;
			29680: outdata = 32'd35856;
			29681: outdata = 32'd35855;
			29682: outdata = 32'd35854;
			29683: outdata = 32'd35853;
			29684: outdata = 32'd35852;
			29685: outdata = 32'd35851;
			29686: outdata = 32'd35850;
			29687: outdata = 32'd35849;
			29688: outdata = 32'd35848;
			29689: outdata = 32'd35847;
			29690: outdata = 32'd35846;
			29691: outdata = 32'd35845;
			29692: outdata = 32'd35844;
			29693: outdata = 32'd35843;
			29694: outdata = 32'd35842;
			29695: outdata = 32'd35841;
			29696: outdata = 32'd35840;
			29697: outdata = 32'd35839;
			29698: outdata = 32'd35838;
			29699: outdata = 32'd35837;
			29700: outdata = 32'd35836;
			29701: outdata = 32'd35835;
			29702: outdata = 32'd35834;
			29703: outdata = 32'd35833;
			29704: outdata = 32'd35832;
			29705: outdata = 32'd35831;
			29706: outdata = 32'd35830;
			29707: outdata = 32'd35829;
			29708: outdata = 32'd35828;
			29709: outdata = 32'd35827;
			29710: outdata = 32'd35826;
			29711: outdata = 32'd35825;
			29712: outdata = 32'd35824;
			29713: outdata = 32'd35823;
			29714: outdata = 32'd35822;
			29715: outdata = 32'd35821;
			29716: outdata = 32'd35820;
			29717: outdata = 32'd35819;
			29718: outdata = 32'd35818;
			29719: outdata = 32'd35817;
			29720: outdata = 32'd35816;
			29721: outdata = 32'd35815;
			29722: outdata = 32'd35814;
			29723: outdata = 32'd35813;
			29724: outdata = 32'd35812;
			29725: outdata = 32'd35811;
			29726: outdata = 32'd35810;
			29727: outdata = 32'd35809;
			29728: outdata = 32'd35808;
			29729: outdata = 32'd35807;
			29730: outdata = 32'd35806;
			29731: outdata = 32'd35805;
			29732: outdata = 32'd35804;
			29733: outdata = 32'd35803;
			29734: outdata = 32'd35802;
			29735: outdata = 32'd35801;
			29736: outdata = 32'd35800;
			29737: outdata = 32'd35799;
			29738: outdata = 32'd35798;
			29739: outdata = 32'd35797;
			29740: outdata = 32'd35796;
			29741: outdata = 32'd35795;
			29742: outdata = 32'd35794;
			29743: outdata = 32'd35793;
			29744: outdata = 32'd35792;
			29745: outdata = 32'd35791;
			29746: outdata = 32'd35790;
			29747: outdata = 32'd35789;
			29748: outdata = 32'd35788;
			29749: outdata = 32'd35787;
			29750: outdata = 32'd35786;
			29751: outdata = 32'd35785;
			29752: outdata = 32'd35784;
			29753: outdata = 32'd35783;
			29754: outdata = 32'd35782;
			29755: outdata = 32'd35781;
			29756: outdata = 32'd35780;
			29757: outdata = 32'd35779;
			29758: outdata = 32'd35778;
			29759: outdata = 32'd35777;
			29760: outdata = 32'd35776;
			29761: outdata = 32'd35775;
			29762: outdata = 32'd35774;
			29763: outdata = 32'd35773;
			29764: outdata = 32'd35772;
			29765: outdata = 32'd35771;
			29766: outdata = 32'd35770;
			29767: outdata = 32'd35769;
			29768: outdata = 32'd35768;
			29769: outdata = 32'd35767;
			29770: outdata = 32'd35766;
			29771: outdata = 32'd35765;
			29772: outdata = 32'd35764;
			29773: outdata = 32'd35763;
			29774: outdata = 32'd35762;
			29775: outdata = 32'd35761;
			29776: outdata = 32'd35760;
			29777: outdata = 32'd35759;
			29778: outdata = 32'd35758;
			29779: outdata = 32'd35757;
			29780: outdata = 32'd35756;
			29781: outdata = 32'd35755;
			29782: outdata = 32'd35754;
			29783: outdata = 32'd35753;
			29784: outdata = 32'd35752;
			29785: outdata = 32'd35751;
			29786: outdata = 32'd35750;
			29787: outdata = 32'd35749;
			29788: outdata = 32'd35748;
			29789: outdata = 32'd35747;
			29790: outdata = 32'd35746;
			29791: outdata = 32'd35745;
			29792: outdata = 32'd35744;
			29793: outdata = 32'd35743;
			29794: outdata = 32'd35742;
			29795: outdata = 32'd35741;
			29796: outdata = 32'd35740;
			29797: outdata = 32'd35739;
			29798: outdata = 32'd35738;
			29799: outdata = 32'd35737;
			29800: outdata = 32'd35736;
			29801: outdata = 32'd35735;
			29802: outdata = 32'd35734;
			29803: outdata = 32'd35733;
			29804: outdata = 32'd35732;
			29805: outdata = 32'd35731;
			29806: outdata = 32'd35730;
			29807: outdata = 32'd35729;
			29808: outdata = 32'd35728;
			29809: outdata = 32'd35727;
			29810: outdata = 32'd35726;
			29811: outdata = 32'd35725;
			29812: outdata = 32'd35724;
			29813: outdata = 32'd35723;
			29814: outdata = 32'd35722;
			29815: outdata = 32'd35721;
			29816: outdata = 32'd35720;
			29817: outdata = 32'd35719;
			29818: outdata = 32'd35718;
			29819: outdata = 32'd35717;
			29820: outdata = 32'd35716;
			29821: outdata = 32'd35715;
			29822: outdata = 32'd35714;
			29823: outdata = 32'd35713;
			29824: outdata = 32'd35712;
			29825: outdata = 32'd35711;
			29826: outdata = 32'd35710;
			29827: outdata = 32'd35709;
			29828: outdata = 32'd35708;
			29829: outdata = 32'd35707;
			29830: outdata = 32'd35706;
			29831: outdata = 32'd35705;
			29832: outdata = 32'd35704;
			29833: outdata = 32'd35703;
			29834: outdata = 32'd35702;
			29835: outdata = 32'd35701;
			29836: outdata = 32'd35700;
			29837: outdata = 32'd35699;
			29838: outdata = 32'd35698;
			29839: outdata = 32'd35697;
			29840: outdata = 32'd35696;
			29841: outdata = 32'd35695;
			29842: outdata = 32'd35694;
			29843: outdata = 32'd35693;
			29844: outdata = 32'd35692;
			29845: outdata = 32'd35691;
			29846: outdata = 32'd35690;
			29847: outdata = 32'd35689;
			29848: outdata = 32'd35688;
			29849: outdata = 32'd35687;
			29850: outdata = 32'd35686;
			29851: outdata = 32'd35685;
			29852: outdata = 32'd35684;
			29853: outdata = 32'd35683;
			29854: outdata = 32'd35682;
			29855: outdata = 32'd35681;
			29856: outdata = 32'd35680;
			29857: outdata = 32'd35679;
			29858: outdata = 32'd35678;
			29859: outdata = 32'd35677;
			29860: outdata = 32'd35676;
			29861: outdata = 32'd35675;
			29862: outdata = 32'd35674;
			29863: outdata = 32'd35673;
			29864: outdata = 32'd35672;
			29865: outdata = 32'd35671;
			29866: outdata = 32'd35670;
			29867: outdata = 32'd35669;
			29868: outdata = 32'd35668;
			29869: outdata = 32'd35667;
			29870: outdata = 32'd35666;
			29871: outdata = 32'd35665;
			29872: outdata = 32'd35664;
			29873: outdata = 32'd35663;
			29874: outdata = 32'd35662;
			29875: outdata = 32'd35661;
			29876: outdata = 32'd35660;
			29877: outdata = 32'd35659;
			29878: outdata = 32'd35658;
			29879: outdata = 32'd35657;
			29880: outdata = 32'd35656;
			29881: outdata = 32'd35655;
			29882: outdata = 32'd35654;
			29883: outdata = 32'd35653;
			29884: outdata = 32'd35652;
			29885: outdata = 32'd35651;
			29886: outdata = 32'd35650;
			29887: outdata = 32'd35649;
			29888: outdata = 32'd35648;
			29889: outdata = 32'd35647;
			29890: outdata = 32'd35646;
			29891: outdata = 32'd35645;
			29892: outdata = 32'd35644;
			29893: outdata = 32'd35643;
			29894: outdata = 32'd35642;
			29895: outdata = 32'd35641;
			29896: outdata = 32'd35640;
			29897: outdata = 32'd35639;
			29898: outdata = 32'd35638;
			29899: outdata = 32'd35637;
			29900: outdata = 32'd35636;
			29901: outdata = 32'd35635;
			29902: outdata = 32'd35634;
			29903: outdata = 32'd35633;
			29904: outdata = 32'd35632;
			29905: outdata = 32'd35631;
			29906: outdata = 32'd35630;
			29907: outdata = 32'd35629;
			29908: outdata = 32'd35628;
			29909: outdata = 32'd35627;
			29910: outdata = 32'd35626;
			29911: outdata = 32'd35625;
			29912: outdata = 32'd35624;
			29913: outdata = 32'd35623;
			29914: outdata = 32'd35622;
			29915: outdata = 32'd35621;
			29916: outdata = 32'd35620;
			29917: outdata = 32'd35619;
			29918: outdata = 32'd35618;
			29919: outdata = 32'd35617;
			29920: outdata = 32'd35616;
			29921: outdata = 32'd35615;
			29922: outdata = 32'd35614;
			29923: outdata = 32'd35613;
			29924: outdata = 32'd35612;
			29925: outdata = 32'd35611;
			29926: outdata = 32'd35610;
			29927: outdata = 32'd35609;
			29928: outdata = 32'd35608;
			29929: outdata = 32'd35607;
			29930: outdata = 32'd35606;
			29931: outdata = 32'd35605;
			29932: outdata = 32'd35604;
			29933: outdata = 32'd35603;
			29934: outdata = 32'd35602;
			29935: outdata = 32'd35601;
			29936: outdata = 32'd35600;
			29937: outdata = 32'd35599;
			29938: outdata = 32'd35598;
			29939: outdata = 32'd35597;
			29940: outdata = 32'd35596;
			29941: outdata = 32'd35595;
			29942: outdata = 32'd35594;
			29943: outdata = 32'd35593;
			29944: outdata = 32'd35592;
			29945: outdata = 32'd35591;
			29946: outdata = 32'd35590;
			29947: outdata = 32'd35589;
			29948: outdata = 32'd35588;
			29949: outdata = 32'd35587;
			29950: outdata = 32'd35586;
			29951: outdata = 32'd35585;
			29952: outdata = 32'd35584;
			29953: outdata = 32'd35583;
			29954: outdata = 32'd35582;
			29955: outdata = 32'd35581;
			29956: outdata = 32'd35580;
			29957: outdata = 32'd35579;
			29958: outdata = 32'd35578;
			29959: outdata = 32'd35577;
			29960: outdata = 32'd35576;
			29961: outdata = 32'd35575;
			29962: outdata = 32'd35574;
			29963: outdata = 32'd35573;
			29964: outdata = 32'd35572;
			29965: outdata = 32'd35571;
			29966: outdata = 32'd35570;
			29967: outdata = 32'd35569;
			29968: outdata = 32'd35568;
			29969: outdata = 32'd35567;
			29970: outdata = 32'd35566;
			29971: outdata = 32'd35565;
			29972: outdata = 32'd35564;
			29973: outdata = 32'd35563;
			29974: outdata = 32'd35562;
			29975: outdata = 32'd35561;
			29976: outdata = 32'd35560;
			29977: outdata = 32'd35559;
			29978: outdata = 32'd35558;
			29979: outdata = 32'd35557;
			29980: outdata = 32'd35556;
			29981: outdata = 32'd35555;
			29982: outdata = 32'd35554;
			29983: outdata = 32'd35553;
			29984: outdata = 32'd35552;
			29985: outdata = 32'd35551;
			29986: outdata = 32'd35550;
			29987: outdata = 32'd35549;
			29988: outdata = 32'd35548;
			29989: outdata = 32'd35547;
			29990: outdata = 32'd35546;
			29991: outdata = 32'd35545;
			29992: outdata = 32'd35544;
			29993: outdata = 32'd35543;
			29994: outdata = 32'd35542;
			29995: outdata = 32'd35541;
			29996: outdata = 32'd35540;
			29997: outdata = 32'd35539;
			29998: outdata = 32'd35538;
			29999: outdata = 32'd35537;
			30000: outdata = 32'd35536;
			30001: outdata = 32'd35535;
			30002: outdata = 32'd35534;
			30003: outdata = 32'd35533;
			30004: outdata = 32'd35532;
			30005: outdata = 32'd35531;
			30006: outdata = 32'd35530;
			30007: outdata = 32'd35529;
			30008: outdata = 32'd35528;
			30009: outdata = 32'd35527;
			30010: outdata = 32'd35526;
			30011: outdata = 32'd35525;
			30012: outdata = 32'd35524;
			30013: outdata = 32'd35523;
			30014: outdata = 32'd35522;
			30015: outdata = 32'd35521;
			30016: outdata = 32'd35520;
			30017: outdata = 32'd35519;
			30018: outdata = 32'd35518;
			30019: outdata = 32'd35517;
			30020: outdata = 32'd35516;
			30021: outdata = 32'd35515;
			30022: outdata = 32'd35514;
			30023: outdata = 32'd35513;
			30024: outdata = 32'd35512;
			30025: outdata = 32'd35511;
			30026: outdata = 32'd35510;
			30027: outdata = 32'd35509;
			30028: outdata = 32'd35508;
			30029: outdata = 32'd35507;
			30030: outdata = 32'd35506;
			30031: outdata = 32'd35505;
			30032: outdata = 32'd35504;
			30033: outdata = 32'd35503;
			30034: outdata = 32'd35502;
			30035: outdata = 32'd35501;
			30036: outdata = 32'd35500;
			30037: outdata = 32'd35499;
			30038: outdata = 32'd35498;
			30039: outdata = 32'd35497;
			30040: outdata = 32'd35496;
			30041: outdata = 32'd35495;
			30042: outdata = 32'd35494;
			30043: outdata = 32'd35493;
			30044: outdata = 32'd35492;
			30045: outdata = 32'd35491;
			30046: outdata = 32'd35490;
			30047: outdata = 32'd35489;
			30048: outdata = 32'd35488;
			30049: outdata = 32'd35487;
			30050: outdata = 32'd35486;
			30051: outdata = 32'd35485;
			30052: outdata = 32'd35484;
			30053: outdata = 32'd35483;
			30054: outdata = 32'd35482;
			30055: outdata = 32'd35481;
			30056: outdata = 32'd35480;
			30057: outdata = 32'd35479;
			30058: outdata = 32'd35478;
			30059: outdata = 32'd35477;
			30060: outdata = 32'd35476;
			30061: outdata = 32'd35475;
			30062: outdata = 32'd35474;
			30063: outdata = 32'd35473;
			30064: outdata = 32'd35472;
			30065: outdata = 32'd35471;
			30066: outdata = 32'd35470;
			30067: outdata = 32'd35469;
			30068: outdata = 32'd35468;
			30069: outdata = 32'd35467;
			30070: outdata = 32'd35466;
			30071: outdata = 32'd35465;
			30072: outdata = 32'd35464;
			30073: outdata = 32'd35463;
			30074: outdata = 32'd35462;
			30075: outdata = 32'd35461;
			30076: outdata = 32'd35460;
			30077: outdata = 32'd35459;
			30078: outdata = 32'd35458;
			30079: outdata = 32'd35457;
			30080: outdata = 32'd35456;
			30081: outdata = 32'd35455;
			30082: outdata = 32'd35454;
			30083: outdata = 32'd35453;
			30084: outdata = 32'd35452;
			30085: outdata = 32'd35451;
			30086: outdata = 32'd35450;
			30087: outdata = 32'd35449;
			30088: outdata = 32'd35448;
			30089: outdata = 32'd35447;
			30090: outdata = 32'd35446;
			30091: outdata = 32'd35445;
			30092: outdata = 32'd35444;
			30093: outdata = 32'd35443;
			30094: outdata = 32'd35442;
			30095: outdata = 32'd35441;
			30096: outdata = 32'd35440;
			30097: outdata = 32'd35439;
			30098: outdata = 32'd35438;
			30099: outdata = 32'd35437;
			30100: outdata = 32'd35436;
			30101: outdata = 32'd35435;
			30102: outdata = 32'd35434;
			30103: outdata = 32'd35433;
			30104: outdata = 32'd35432;
			30105: outdata = 32'd35431;
			30106: outdata = 32'd35430;
			30107: outdata = 32'd35429;
			30108: outdata = 32'd35428;
			30109: outdata = 32'd35427;
			30110: outdata = 32'd35426;
			30111: outdata = 32'd35425;
			30112: outdata = 32'd35424;
			30113: outdata = 32'd35423;
			30114: outdata = 32'd35422;
			30115: outdata = 32'd35421;
			30116: outdata = 32'd35420;
			30117: outdata = 32'd35419;
			30118: outdata = 32'd35418;
			30119: outdata = 32'd35417;
			30120: outdata = 32'd35416;
			30121: outdata = 32'd35415;
			30122: outdata = 32'd35414;
			30123: outdata = 32'd35413;
			30124: outdata = 32'd35412;
			30125: outdata = 32'd35411;
			30126: outdata = 32'd35410;
			30127: outdata = 32'd35409;
			30128: outdata = 32'd35408;
			30129: outdata = 32'd35407;
			30130: outdata = 32'd35406;
			30131: outdata = 32'd35405;
			30132: outdata = 32'd35404;
			30133: outdata = 32'd35403;
			30134: outdata = 32'd35402;
			30135: outdata = 32'd35401;
			30136: outdata = 32'd35400;
			30137: outdata = 32'd35399;
			30138: outdata = 32'd35398;
			30139: outdata = 32'd35397;
			30140: outdata = 32'd35396;
			30141: outdata = 32'd35395;
			30142: outdata = 32'd35394;
			30143: outdata = 32'd35393;
			30144: outdata = 32'd35392;
			30145: outdata = 32'd35391;
			30146: outdata = 32'd35390;
			30147: outdata = 32'd35389;
			30148: outdata = 32'd35388;
			30149: outdata = 32'd35387;
			30150: outdata = 32'd35386;
			30151: outdata = 32'd35385;
			30152: outdata = 32'd35384;
			30153: outdata = 32'd35383;
			30154: outdata = 32'd35382;
			30155: outdata = 32'd35381;
			30156: outdata = 32'd35380;
			30157: outdata = 32'd35379;
			30158: outdata = 32'd35378;
			30159: outdata = 32'd35377;
			30160: outdata = 32'd35376;
			30161: outdata = 32'd35375;
			30162: outdata = 32'd35374;
			30163: outdata = 32'd35373;
			30164: outdata = 32'd35372;
			30165: outdata = 32'd35371;
			30166: outdata = 32'd35370;
			30167: outdata = 32'd35369;
			30168: outdata = 32'd35368;
			30169: outdata = 32'd35367;
			30170: outdata = 32'd35366;
			30171: outdata = 32'd35365;
			30172: outdata = 32'd35364;
			30173: outdata = 32'd35363;
			30174: outdata = 32'd35362;
			30175: outdata = 32'd35361;
			30176: outdata = 32'd35360;
			30177: outdata = 32'd35359;
			30178: outdata = 32'd35358;
			30179: outdata = 32'd35357;
			30180: outdata = 32'd35356;
			30181: outdata = 32'd35355;
			30182: outdata = 32'd35354;
			30183: outdata = 32'd35353;
			30184: outdata = 32'd35352;
			30185: outdata = 32'd35351;
			30186: outdata = 32'd35350;
			30187: outdata = 32'd35349;
			30188: outdata = 32'd35348;
			30189: outdata = 32'd35347;
			30190: outdata = 32'd35346;
			30191: outdata = 32'd35345;
			30192: outdata = 32'd35344;
			30193: outdata = 32'd35343;
			30194: outdata = 32'd35342;
			30195: outdata = 32'd35341;
			30196: outdata = 32'd35340;
			30197: outdata = 32'd35339;
			30198: outdata = 32'd35338;
			30199: outdata = 32'd35337;
			30200: outdata = 32'd35336;
			30201: outdata = 32'd35335;
			30202: outdata = 32'd35334;
			30203: outdata = 32'd35333;
			30204: outdata = 32'd35332;
			30205: outdata = 32'd35331;
			30206: outdata = 32'd35330;
			30207: outdata = 32'd35329;
			30208: outdata = 32'd35328;
			30209: outdata = 32'd35327;
			30210: outdata = 32'd35326;
			30211: outdata = 32'd35325;
			30212: outdata = 32'd35324;
			30213: outdata = 32'd35323;
			30214: outdata = 32'd35322;
			30215: outdata = 32'd35321;
			30216: outdata = 32'd35320;
			30217: outdata = 32'd35319;
			30218: outdata = 32'd35318;
			30219: outdata = 32'd35317;
			30220: outdata = 32'd35316;
			30221: outdata = 32'd35315;
			30222: outdata = 32'd35314;
			30223: outdata = 32'd35313;
			30224: outdata = 32'd35312;
			30225: outdata = 32'd35311;
			30226: outdata = 32'd35310;
			30227: outdata = 32'd35309;
			30228: outdata = 32'd35308;
			30229: outdata = 32'd35307;
			30230: outdata = 32'd35306;
			30231: outdata = 32'd35305;
			30232: outdata = 32'd35304;
			30233: outdata = 32'd35303;
			30234: outdata = 32'd35302;
			30235: outdata = 32'd35301;
			30236: outdata = 32'd35300;
			30237: outdata = 32'd35299;
			30238: outdata = 32'd35298;
			30239: outdata = 32'd35297;
			30240: outdata = 32'd35296;
			30241: outdata = 32'd35295;
			30242: outdata = 32'd35294;
			30243: outdata = 32'd35293;
			30244: outdata = 32'd35292;
			30245: outdata = 32'd35291;
			30246: outdata = 32'd35290;
			30247: outdata = 32'd35289;
			30248: outdata = 32'd35288;
			30249: outdata = 32'd35287;
			30250: outdata = 32'd35286;
			30251: outdata = 32'd35285;
			30252: outdata = 32'd35284;
			30253: outdata = 32'd35283;
			30254: outdata = 32'd35282;
			30255: outdata = 32'd35281;
			30256: outdata = 32'd35280;
			30257: outdata = 32'd35279;
			30258: outdata = 32'd35278;
			30259: outdata = 32'd35277;
			30260: outdata = 32'd35276;
			30261: outdata = 32'd35275;
			30262: outdata = 32'd35274;
			30263: outdata = 32'd35273;
			30264: outdata = 32'd35272;
			30265: outdata = 32'd35271;
			30266: outdata = 32'd35270;
			30267: outdata = 32'd35269;
			30268: outdata = 32'd35268;
			30269: outdata = 32'd35267;
			30270: outdata = 32'd35266;
			30271: outdata = 32'd35265;
			30272: outdata = 32'd35264;
			30273: outdata = 32'd35263;
			30274: outdata = 32'd35262;
			30275: outdata = 32'd35261;
			30276: outdata = 32'd35260;
			30277: outdata = 32'd35259;
			30278: outdata = 32'd35258;
			30279: outdata = 32'd35257;
			30280: outdata = 32'd35256;
			30281: outdata = 32'd35255;
			30282: outdata = 32'd35254;
			30283: outdata = 32'd35253;
			30284: outdata = 32'd35252;
			30285: outdata = 32'd35251;
			30286: outdata = 32'd35250;
			30287: outdata = 32'd35249;
			30288: outdata = 32'd35248;
			30289: outdata = 32'd35247;
			30290: outdata = 32'd35246;
			30291: outdata = 32'd35245;
			30292: outdata = 32'd35244;
			30293: outdata = 32'd35243;
			30294: outdata = 32'd35242;
			30295: outdata = 32'd35241;
			30296: outdata = 32'd35240;
			30297: outdata = 32'd35239;
			30298: outdata = 32'd35238;
			30299: outdata = 32'd35237;
			30300: outdata = 32'd35236;
			30301: outdata = 32'd35235;
			30302: outdata = 32'd35234;
			30303: outdata = 32'd35233;
			30304: outdata = 32'd35232;
			30305: outdata = 32'd35231;
			30306: outdata = 32'd35230;
			30307: outdata = 32'd35229;
			30308: outdata = 32'd35228;
			30309: outdata = 32'd35227;
			30310: outdata = 32'd35226;
			30311: outdata = 32'd35225;
			30312: outdata = 32'd35224;
			30313: outdata = 32'd35223;
			30314: outdata = 32'd35222;
			30315: outdata = 32'd35221;
			30316: outdata = 32'd35220;
			30317: outdata = 32'd35219;
			30318: outdata = 32'd35218;
			30319: outdata = 32'd35217;
			30320: outdata = 32'd35216;
			30321: outdata = 32'd35215;
			30322: outdata = 32'd35214;
			30323: outdata = 32'd35213;
			30324: outdata = 32'd35212;
			30325: outdata = 32'd35211;
			30326: outdata = 32'd35210;
			30327: outdata = 32'd35209;
			30328: outdata = 32'd35208;
			30329: outdata = 32'd35207;
			30330: outdata = 32'd35206;
			30331: outdata = 32'd35205;
			30332: outdata = 32'd35204;
			30333: outdata = 32'd35203;
			30334: outdata = 32'd35202;
			30335: outdata = 32'd35201;
			30336: outdata = 32'd35200;
			30337: outdata = 32'd35199;
			30338: outdata = 32'd35198;
			30339: outdata = 32'd35197;
			30340: outdata = 32'd35196;
			30341: outdata = 32'd35195;
			30342: outdata = 32'd35194;
			30343: outdata = 32'd35193;
			30344: outdata = 32'd35192;
			30345: outdata = 32'd35191;
			30346: outdata = 32'd35190;
			30347: outdata = 32'd35189;
			30348: outdata = 32'd35188;
			30349: outdata = 32'd35187;
			30350: outdata = 32'd35186;
			30351: outdata = 32'd35185;
			30352: outdata = 32'd35184;
			30353: outdata = 32'd35183;
			30354: outdata = 32'd35182;
			30355: outdata = 32'd35181;
			30356: outdata = 32'd35180;
			30357: outdata = 32'd35179;
			30358: outdata = 32'd35178;
			30359: outdata = 32'd35177;
			30360: outdata = 32'd35176;
			30361: outdata = 32'd35175;
			30362: outdata = 32'd35174;
			30363: outdata = 32'd35173;
			30364: outdata = 32'd35172;
			30365: outdata = 32'd35171;
			30366: outdata = 32'd35170;
			30367: outdata = 32'd35169;
			30368: outdata = 32'd35168;
			30369: outdata = 32'd35167;
			30370: outdata = 32'd35166;
			30371: outdata = 32'd35165;
			30372: outdata = 32'd35164;
			30373: outdata = 32'd35163;
			30374: outdata = 32'd35162;
			30375: outdata = 32'd35161;
			30376: outdata = 32'd35160;
			30377: outdata = 32'd35159;
			30378: outdata = 32'd35158;
			30379: outdata = 32'd35157;
			30380: outdata = 32'd35156;
			30381: outdata = 32'd35155;
			30382: outdata = 32'd35154;
			30383: outdata = 32'd35153;
			30384: outdata = 32'd35152;
			30385: outdata = 32'd35151;
			30386: outdata = 32'd35150;
			30387: outdata = 32'd35149;
			30388: outdata = 32'd35148;
			30389: outdata = 32'd35147;
			30390: outdata = 32'd35146;
			30391: outdata = 32'd35145;
			30392: outdata = 32'd35144;
			30393: outdata = 32'd35143;
			30394: outdata = 32'd35142;
			30395: outdata = 32'd35141;
			30396: outdata = 32'd35140;
			30397: outdata = 32'd35139;
			30398: outdata = 32'd35138;
			30399: outdata = 32'd35137;
			30400: outdata = 32'd35136;
			30401: outdata = 32'd35135;
			30402: outdata = 32'd35134;
			30403: outdata = 32'd35133;
			30404: outdata = 32'd35132;
			30405: outdata = 32'd35131;
			30406: outdata = 32'd35130;
			30407: outdata = 32'd35129;
			30408: outdata = 32'd35128;
			30409: outdata = 32'd35127;
			30410: outdata = 32'd35126;
			30411: outdata = 32'd35125;
			30412: outdata = 32'd35124;
			30413: outdata = 32'd35123;
			30414: outdata = 32'd35122;
			30415: outdata = 32'd35121;
			30416: outdata = 32'd35120;
			30417: outdata = 32'd35119;
			30418: outdata = 32'd35118;
			30419: outdata = 32'd35117;
			30420: outdata = 32'd35116;
			30421: outdata = 32'd35115;
			30422: outdata = 32'd35114;
			30423: outdata = 32'd35113;
			30424: outdata = 32'd35112;
			30425: outdata = 32'd35111;
			30426: outdata = 32'd35110;
			30427: outdata = 32'd35109;
			30428: outdata = 32'd35108;
			30429: outdata = 32'd35107;
			30430: outdata = 32'd35106;
			30431: outdata = 32'd35105;
			30432: outdata = 32'd35104;
			30433: outdata = 32'd35103;
			30434: outdata = 32'd35102;
			30435: outdata = 32'd35101;
			30436: outdata = 32'd35100;
			30437: outdata = 32'd35099;
			30438: outdata = 32'd35098;
			30439: outdata = 32'd35097;
			30440: outdata = 32'd35096;
			30441: outdata = 32'd35095;
			30442: outdata = 32'd35094;
			30443: outdata = 32'd35093;
			30444: outdata = 32'd35092;
			30445: outdata = 32'd35091;
			30446: outdata = 32'd35090;
			30447: outdata = 32'd35089;
			30448: outdata = 32'd35088;
			30449: outdata = 32'd35087;
			30450: outdata = 32'd35086;
			30451: outdata = 32'd35085;
			30452: outdata = 32'd35084;
			30453: outdata = 32'd35083;
			30454: outdata = 32'd35082;
			30455: outdata = 32'd35081;
			30456: outdata = 32'd35080;
			30457: outdata = 32'd35079;
			30458: outdata = 32'd35078;
			30459: outdata = 32'd35077;
			30460: outdata = 32'd35076;
			30461: outdata = 32'd35075;
			30462: outdata = 32'd35074;
			30463: outdata = 32'd35073;
			30464: outdata = 32'd35072;
			30465: outdata = 32'd35071;
			30466: outdata = 32'd35070;
			30467: outdata = 32'd35069;
			30468: outdata = 32'd35068;
			30469: outdata = 32'd35067;
			30470: outdata = 32'd35066;
			30471: outdata = 32'd35065;
			30472: outdata = 32'd35064;
			30473: outdata = 32'd35063;
			30474: outdata = 32'd35062;
			30475: outdata = 32'd35061;
			30476: outdata = 32'd35060;
			30477: outdata = 32'd35059;
			30478: outdata = 32'd35058;
			30479: outdata = 32'd35057;
			30480: outdata = 32'd35056;
			30481: outdata = 32'd35055;
			30482: outdata = 32'd35054;
			30483: outdata = 32'd35053;
			30484: outdata = 32'd35052;
			30485: outdata = 32'd35051;
			30486: outdata = 32'd35050;
			30487: outdata = 32'd35049;
			30488: outdata = 32'd35048;
			30489: outdata = 32'd35047;
			30490: outdata = 32'd35046;
			30491: outdata = 32'd35045;
			30492: outdata = 32'd35044;
			30493: outdata = 32'd35043;
			30494: outdata = 32'd35042;
			30495: outdata = 32'd35041;
			30496: outdata = 32'd35040;
			30497: outdata = 32'd35039;
			30498: outdata = 32'd35038;
			30499: outdata = 32'd35037;
			30500: outdata = 32'd35036;
			30501: outdata = 32'd35035;
			30502: outdata = 32'd35034;
			30503: outdata = 32'd35033;
			30504: outdata = 32'd35032;
			30505: outdata = 32'd35031;
			30506: outdata = 32'd35030;
			30507: outdata = 32'd35029;
			30508: outdata = 32'd35028;
			30509: outdata = 32'd35027;
			30510: outdata = 32'd35026;
			30511: outdata = 32'd35025;
			30512: outdata = 32'd35024;
			30513: outdata = 32'd35023;
			30514: outdata = 32'd35022;
			30515: outdata = 32'd35021;
			30516: outdata = 32'd35020;
			30517: outdata = 32'd35019;
			30518: outdata = 32'd35018;
			30519: outdata = 32'd35017;
			30520: outdata = 32'd35016;
			30521: outdata = 32'd35015;
			30522: outdata = 32'd35014;
			30523: outdata = 32'd35013;
			30524: outdata = 32'd35012;
			30525: outdata = 32'd35011;
			30526: outdata = 32'd35010;
			30527: outdata = 32'd35009;
			30528: outdata = 32'd35008;
			30529: outdata = 32'd35007;
			30530: outdata = 32'd35006;
			30531: outdata = 32'd35005;
			30532: outdata = 32'd35004;
			30533: outdata = 32'd35003;
			30534: outdata = 32'd35002;
			30535: outdata = 32'd35001;
			30536: outdata = 32'd35000;
			30537: outdata = 32'd34999;
			30538: outdata = 32'd34998;
			30539: outdata = 32'd34997;
			30540: outdata = 32'd34996;
			30541: outdata = 32'd34995;
			30542: outdata = 32'd34994;
			30543: outdata = 32'd34993;
			30544: outdata = 32'd34992;
			30545: outdata = 32'd34991;
			30546: outdata = 32'd34990;
			30547: outdata = 32'd34989;
			30548: outdata = 32'd34988;
			30549: outdata = 32'd34987;
			30550: outdata = 32'd34986;
			30551: outdata = 32'd34985;
			30552: outdata = 32'd34984;
			30553: outdata = 32'd34983;
			30554: outdata = 32'd34982;
			30555: outdata = 32'd34981;
			30556: outdata = 32'd34980;
			30557: outdata = 32'd34979;
			30558: outdata = 32'd34978;
			30559: outdata = 32'd34977;
			30560: outdata = 32'd34976;
			30561: outdata = 32'd34975;
			30562: outdata = 32'd34974;
			30563: outdata = 32'd34973;
			30564: outdata = 32'd34972;
			30565: outdata = 32'd34971;
			30566: outdata = 32'd34970;
			30567: outdata = 32'd34969;
			30568: outdata = 32'd34968;
			30569: outdata = 32'd34967;
			30570: outdata = 32'd34966;
			30571: outdata = 32'd34965;
			30572: outdata = 32'd34964;
			30573: outdata = 32'd34963;
			30574: outdata = 32'd34962;
			30575: outdata = 32'd34961;
			30576: outdata = 32'd34960;
			30577: outdata = 32'd34959;
			30578: outdata = 32'd34958;
			30579: outdata = 32'd34957;
			30580: outdata = 32'd34956;
			30581: outdata = 32'd34955;
			30582: outdata = 32'd34954;
			30583: outdata = 32'd34953;
			30584: outdata = 32'd34952;
			30585: outdata = 32'd34951;
			30586: outdata = 32'd34950;
			30587: outdata = 32'd34949;
			30588: outdata = 32'd34948;
			30589: outdata = 32'd34947;
			30590: outdata = 32'd34946;
			30591: outdata = 32'd34945;
			30592: outdata = 32'd34944;
			30593: outdata = 32'd34943;
			30594: outdata = 32'd34942;
			30595: outdata = 32'd34941;
			30596: outdata = 32'd34940;
			30597: outdata = 32'd34939;
			30598: outdata = 32'd34938;
			30599: outdata = 32'd34937;
			30600: outdata = 32'd34936;
			30601: outdata = 32'd34935;
			30602: outdata = 32'd34934;
			30603: outdata = 32'd34933;
			30604: outdata = 32'd34932;
			30605: outdata = 32'd34931;
			30606: outdata = 32'd34930;
			30607: outdata = 32'd34929;
			30608: outdata = 32'd34928;
			30609: outdata = 32'd34927;
			30610: outdata = 32'd34926;
			30611: outdata = 32'd34925;
			30612: outdata = 32'd34924;
			30613: outdata = 32'd34923;
			30614: outdata = 32'd34922;
			30615: outdata = 32'd34921;
			30616: outdata = 32'd34920;
			30617: outdata = 32'd34919;
			30618: outdata = 32'd34918;
			30619: outdata = 32'd34917;
			30620: outdata = 32'd34916;
			30621: outdata = 32'd34915;
			30622: outdata = 32'd34914;
			30623: outdata = 32'd34913;
			30624: outdata = 32'd34912;
			30625: outdata = 32'd34911;
			30626: outdata = 32'd34910;
			30627: outdata = 32'd34909;
			30628: outdata = 32'd34908;
			30629: outdata = 32'd34907;
			30630: outdata = 32'd34906;
			30631: outdata = 32'd34905;
			30632: outdata = 32'd34904;
			30633: outdata = 32'd34903;
			30634: outdata = 32'd34902;
			30635: outdata = 32'd34901;
			30636: outdata = 32'd34900;
			30637: outdata = 32'd34899;
			30638: outdata = 32'd34898;
			30639: outdata = 32'd34897;
			30640: outdata = 32'd34896;
			30641: outdata = 32'd34895;
			30642: outdata = 32'd34894;
			30643: outdata = 32'd34893;
			30644: outdata = 32'd34892;
			30645: outdata = 32'd34891;
			30646: outdata = 32'd34890;
			30647: outdata = 32'd34889;
			30648: outdata = 32'd34888;
			30649: outdata = 32'd34887;
			30650: outdata = 32'd34886;
			30651: outdata = 32'd34885;
			30652: outdata = 32'd34884;
			30653: outdata = 32'd34883;
			30654: outdata = 32'd34882;
			30655: outdata = 32'd34881;
			30656: outdata = 32'd34880;
			30657: outdata = 32'd34879;
			30658: outdata = 32'd34878;
			30659: outdata = 32'd34877;
			30660: outdata = 32'd34876;
			30661: outdata = 32'd34875;
			30662: outdata = 32'd34874;
			30663: outdata = 32'd34873;
			30664: outdata = 32'd34872;
			30665: outdata = 32'd34871;
			30666: outdata = 32'd34870;
			30667: outdata = 32'd34869;
			30668: outdata = 32'd34868;
			30669: outdata = 32'd34867;
			30670: outdata = 32'd34866;
			30671: outdata = 32'd34865;
			30672: outdata = 32'd34864;
			30673: outdata = 32'd34863;
			30674: outdata = 32'd34862;
			30675: outdata = 32'd34861;
			30676: outdata = 32'd34860;
			30677: outdata = 32'd34859;
			30678: outdata = 32'd34858;
			30679: outdata = 32'd34857;
			30680: outdata = 32'd34856;
			30681: outdata = 32'd34855;
			30682: outdata = 32'd34854;
			30683: outdata = 32'd34853;
			30684: outdata = 32'd34852;
			30685: outdata = 32'd34851;
			30686: outdata = 32'd34850;
			30687: outdata = 32'd34849;
			30688: outdata = 32'd34848;
			30689: outdata = 32'd34847;
			30690: outdata = 32'd34846;
			30691: outdata = 32'd34845;
			30692: outdata = 32'd34844;
			30693: outdata = 32'd34843;
			30694: outdata = 32'd34842;
			30695: outdata = 32'd34841;
			30696: outdata = 32'd34840;
			30697: outdata = 32'd34839;
			30698: outdata = 32'd34838;
			30699: outdata = 32'd34837;
			30700: outdata = 32'd34836;
			30701: outdata = 32'd34835;
			30702: outdata = 32'd34834;
			30703: outdata = 32'd34833;
			30704: outdata = 32'd34832;
			30705: outdata = 32'd34831;
			30706: outdata = 32'd34830;
			30707: outdata = 32'd34829;
			30708: outdata = 32'd34828;
			30709: outdata = 32'd34827;
			30710: outdata = 32'd34826;
			30711: outdata = 32'd34825;
			30712: outdata = 32'd34824;
			30713: outdata = 32'd34823;
			30714: outdata = 32'd34822;
			30715: outdata = 32'd34821;
			30716: outdata = 32'd34820;
			30717: outdata = 32'd34819;
			30718: outdata = 32'd34818;
			30719: outdata = 32'd34817;
			30720: outdata = 32'd34816;
			30721: outdata = 32'd34815;
			30722: outdata = 32'd34814;
			30723: outdata = 32'd34813;
			30724: outdata = 32'd34812;
			30725: outdata = 32'd34811;
			30726: outdata = 32'd34810;
			30727: outdata = 32'd34809;
			30728: outdata = 32'd34808;
			30729: outdata = 32'd34807;
			30730: outdata = 32'd34806;
			30731: outdata = 32'd34805;
			30732: outdata = 32'd34804;
			30733: outdata = 32'd34803;
			30734: outdata = 32'd34802;
			30735: outdata = 32'd34801;
			30736: outdata = 32'd34800;
			30737: outdata = 32'd34799;
			30738: outdata = 32'd34798;
			30739: outdata = 32'd34797;
			30740: outdata = 32'd34796;
			30741: outdata = 32'd34795;
			30742: outdata = 32'd34794;
			30743: outdata = 32'd34793;
			30744: outdata = 32'd34792;
			30745: outdata = 32'd34791;
			30746: outdata = 32'd34790;
			30747: outdata = 32'd34789;
			30748: outdata = 32'd34788;
			30749: outdata = 32'd34787;
			30750: outdata = 32'd34786;
			30751: outdata = 32'd34785;
			30752: outdata = 32'd34784;
			30753: outdata = 32'd34783;
			30754: outdata = 32'd34782;
			30755: outdata = 32'd34781;
			30756: outdata = 32'd34780;
			30757: outdata = 32'd34779;
			30758: outdata = 32'd34778;
			30759: outdata = 32'd34777;
			30760: outdata = 32'd34776;
			30761: outdata = 32'd34775;
			30762: outdata = 32'd34774;
			30763: outdata = 32'd34773;
			30764: outdata = 32'd34772;
			30765: outdata = 32'd34771;
			30766: outdata = 32'd34770;
			30767: outdata = 32'd34769;
			30768: outdata = 32'd34768;
			30769: outdata = 32'd34767;
			30770: outdata = 32'd34766;
			30771: outdata = 32'd34765;
			30772: outdata = 32'd34764;
			30773: outdata = 32'd34763;
			30774: outdata = 32'd34762;
			30775: outdata = 32'd34761;
			30776: outdata = 32'd34760;
			30777: outdata = 32'd34759;
			30778: outdata = 32'd34758;
			30779: outdata = 32'd34757;
			30780: outdata = 32'd34756;
			30781: outdata = 32'd34755;
			30782: outdata = 32'd34754;
			30783: outdata = 32'd34753;
			30784: outdata = 32'd34752;
			30785: outdata = 32'd34751;
			30786: outdata = 32'd34750;
			30787: outdata = 32'd34749;
			30788: outdata = 32'd34748;
			30789: outdata = 32'd34747;
			30790: outdata = 32'd34746;
			30791: outdata = 32'd34745;
			30792: outdata = 32'd34744;
			30793: outdata = 32'd34743;
			30794: outdata = 32'd34742;
			30795: outdata = 32'd34741;
			30796: outdata = 32'd34740;
			30797: outdata = 32'd34739;
			30798: outdata = 32'd34738;
			30799: outdata = 32'd34737;
			30800: outdata = 32'd34736;
			30801: outdata = 32'd34735;
			30802: outdata = 32'd34734;
			30803: outdata = 32'd34733;
			30804: outdata = 32'd34732;
			30805: outdata = 32'd34731;
			30806: outdata = 32'd34730;
			30807: outdata = 32'd34729;
			30808: outdata = 32'd34728;
			30809: outdata = 32'd34727;
			30810: outdata = 32'd34726;
			30811: outdata = 32'd34725;
			30812: outdata = 32'd34724;
			30813: outdata = 32'd34723;
			30814: outdata = 32'd34722;
			30815: outdata = 32'd34721;
			30816: outdata = 32'd34720;
			30817: outdata = 32'd34719;
			30818: outdata = 32'd34718;
			30819: outdata = 32'd34717;
			30820: outdata = 32'd34716;
			30821: outdata = 32'd34715;
			30822: outdata = 32'd34714;
			30823: outdata = 32'd34713;
			30824: outdata = 32'd34712;
			30825: outdata = 32'd34711;
			30826: outdata = 32'd34710;
			30827: outdata = 32'd34709;
			30828: outdata = 32'd34708;
			30829: outdata = 32'd34707;
			30830: outdata = 32'd34706;
			30831: outdata = 32'd34705;
			30832: outdata = 32'd34704;
			30833: outdata = 32'd34703;
			30834: outdata = 32'd34702;
			30835: outdata = 32'd34701;
			30836: outdata = 32'd34700;
			30837: outdata = 32'd34699;
			30838: outdata = 32'd34698;
			30839: outdata = 32'd34697;
			30840: outdata = 32'd34696;
			30841: outdata = 32'd34695;
			30842: outdata = 32'd34694;
			30843: outdata = 32'd34693;
			30844: outdata = 32'd34692;
			30845: outdata = 32'd34691;
			30846: outdata = 32'd34690;
			30847: outdata = 32'd34689;
			30848: outdata = 32'd34688;
			30849: outdata = 32'd34687;
			30850: outdata = 32'd34686;
			30851: outdata = 32'd34685;
			30852: outdata = 32'd34684;
			30853: outdata = 32'd34683;
			30854: outdata = 32'd34682;
			30855: outdata = 32'd34681;
			30856: outdata = 32'd34680;
			30857: outdata = 32'd34679;
			30858: outdata = 32'd34678;
			30859: outdata = 32'd34677;
			30860: outdata = 32'd34676;
			30861: outdata = 32'd34675;
			30862: outdata = 32'd34674;
			30863: outdata = 32'd34673;
			30864: outdata = 32'd34672;
			30865: outdata = 32'd34671;
			30866: outdata = 32'd34670;
			30867: outdata = 32'd34669;
			30868: outdata = 32'd34668;
			30869: outdata = 32'd34667;
			30870: outdata = 32'd34666;
			30871: outdata = 32'd34665;
			30872: outdata = 32'd34664;
			30873: outdata = 32'd34663;
			30874: outdata = 32'd34662;
			30875: outdata = 32'd34661;
			30876: outdata = 32'd34660;
			30877: outdata = 32'd34659;
			30878: outdata = 32'd34658;
			30879: outdata = 32'd34657;
			30880: outdata = 32'd34656;
			30881: outdata = 32'd34655;
			30882: outdata = 32'd34654;
			30883: outdata = 32'd34653;
			30884: outdata = 32'd34652;
			30885: outdata = 32'd34651;
			30886: outdata = 32'd34650;
			30887: outdata = 32'd34649;
			30888: outdata = 32'd34648;
			30889: outdata = 32'd34647;
			30890: outdata = 32'd34646;
			30891: outdata = 32'd34645;
			30892: outdata = 32'd34644;
			30893: outdata = 32'd34643;
			30894: outdata = 32'd34642;
			30895: outdata = 32'd34641;
			30896: outdata = 32'd34640;
			30897: outdata = 32'd34639;
			30898: outdata = 32'd34638;
			30899: outdata = 32'd34637;
			30900: outdata = 32'd34636;
			30901: outdata = 32'd34635;
			30902: outdata = 32'd34634;
			30903: outdata = 32'd34633;
			30904: outdata = 32'd34632;
			30905: outdata = 32'd34631;
			30906: outdata = 32'd34630;
			30907: outdata = 32'd34629;
			30908: outdata = 32'd34628;
			30909: outdata = 32'd34627;
			30910: outdata = 32'd34626;
			30911: outdata = 32'd34625;
			30912: outdata = 32'd34624;
			30913: outdata = 32'd34623;
			30914: outdata = 32'd34622;
			30915: outdata = 32'd34621;
			30916: outdata = 32'd34620;
			30917: outdata = 32'd34619;
			30918: outdata = 32'd34618;
			30919: outdata = 32'd34617;
			30920: outdata = 32'd34616;
			30921: outdata = 32'd34615;
			30922: outdata = 32'd34614;
			30923: outdata = 32'd34613;
			30924: outdata = 32'd34612;
			30925: outdata = 32'd34611;
			30926: outdata = 32'd34610;
			30927: outdata = 32'd34609;
			30928: outdata = 32'd34608;
			30929: outdata = 32'd34607;
			30930: outdata = 32'd34606;
			30931: outdata = 32'd34605;
			30932: outdata = 32'd34604;
			30933: outdata = 32'd34603;
			30934: outdata = 32'd34602;
			30935: outdata = 32'd34601;
			30936: outdata = 32'd34600;
			30937: outdata = 32'd34599;
			30938: outdata = 32'd34598;
			30939: outdata = 32'd34597;
			30940: outdata = 32'd34596;
			30941: outdata = 32'd34595;
			30942: outdata = 32'd34594;
			30943: outdata = 32'd34593;
			30944: outdata = 32'd34592;
			30945: outdata = 32'd34591;
			30946: outdata = 32'd34590;
			30947: outdata = 32'd34589;
			30948: outdata = 32'd34588;
			30949: outdata = 32'd34587;
			30950: outdata = 32'd34586;
			30951: outdata = 32'd34585;
			30952: outdata = 32'd34584;
			30953: outdata = 32'd34583;
			30954: outdata = 32'd34582;
			30955: outdata = 32'd34581;
			30956: outdata = 32'd34580;
			30957: outdata = 32'd34579;
			30958: outdata = 32'd34578;
			30959: outdata = 32'd34577;
			30960: outdata = 32'd34576;
			30961: outdata = 32'd34575;
			30962: outdata = 32'd34574;
			30963: outdata = 32'd34573;
			30964: outdata = 32'd34572;
			30965: outdata = 32'd34571;
			30966: outdata = 32'd34570;
			30967: outdata = 32'd34569;
			30968: outdata = 32'd34568;
			30969: outdata = 32'd34567;
			30970: outdata = 32'd34566;
			30971: outdata = 32'd34565;
			30972: outdata = 32'd34564;
			30973: outdata = 32'd34563;
			30974: outdata = 32'd34562;
			30975: outdata = 32'd34561;
			30976: outdata = 32'd34560;
			30977: outdata = 32'd34559;
			30978: outdata = 32'd34558;
			30979: outdata = 32'd34557;
			30980: outdata = 32'd34556;
			30981: outdata = 32'd34555;
			30982: outdata = 32'd34554;
			30983: outdata = 32'd34553;
			30984: outdata = 32'd34552;
			30985: outdata = 32'd34551;
			30986: outdata = 32'd34550;
			30987: outdata = 32'd34549;
			30988: outdata = 32'd34548;
			30989: outdata = 32'd34547;
			30990: outdata = 32'd34546;
			30991: outdata = 32'd34545;
			30992: outdata = 32'd34544;
			30993: outdata = 32'd34543;
			30994: outdata = 32'd34542;
			30995: outdata = 32'd34541;
			30996: outdata = 32'd34540;
			30997: outdata = 32'd34539;
			30998: outdata = 32'd34538;
			30999: outdata = 32'd34537;
			31000: outdata = 32'd34536;
			31001: outdata = 32'd34535;
			31002: outdata = 32'd34534;
			31003: outdata = 32'd34533;
			31004: outdata = 32'd34532;
			31005: outdata = 32'd34531;
			31006: outdata = 32'd34530;
			31007: outdata = 32'd34529;
			31008: outdata = 32'd34528;
			31009: outdata = 32'd34527;
			31010: outdata = 32'd34526;
			31011: outdata = 32'd34525;
			31012: outdata = 32'd34524;
			31013: outdata = 32'd34523;
			31014: outdata = 32'd34522;
			31015: outdata = 32'd34521;
			31016: outdata = 32'd34520;
			31017: outdata = 32'd34519;
			31018: outdata = 32'd34518;
			31019: outdata = 32'd34517;
			31020: outdata = 32'd34516;
			31021: outdata = 32'd34515;
			31022: outdata = 32'd34514;
			31023: outdata = 32'd34513;
			31024: outdata = 32'd34512;
			31025: outdata = 32'd34511;
			31026: outdata = 32'd34510;
			31027: outdata = 32'd34509;
			31028: outdata = 32'd34508;
			31029: outdata = 32'd34507;
			31030: outdata = 32'd34506;
			31031: outdata = 32'd34505;
			31032: outdata = 32'd34504;
			31033: outdata = 32'd34503;
			31034: outdata = 32'd34502;
			31035: outdata = 32'd34501;
			31036: outdata = 32'd34500;
			31037: outdata = 32'd34499;
			31038: outdata = 32'd34498;
			31039: outdata = 32'd34497;
			31040: outdata = 32'd34496;
			31041: outdata = 32'd34495;
			31042: outdata = 32'd34494;
			31043: outdata = 32'd34493;
			31044: outdata = 32'd34492;
			31045: outdata = 32'd34491;
			31046: outdata = 32'd34490;
			31047: outdata = 32'd34489;
			31048: outdata = 32'd34488;
			31049: outdata = 32'd34487;
			31050: outdata = 32'd34486;
			31051: outdata = 32'd34485;
			31052: outdata = 32'd34484;
			31053: outdata = 32'd34483;
			31054: outdata = 32'd34482;
			31055: outdata = 32'd34481;
			31056: outdata = 32'd34480;
			31057: outdata = 32'd34479;
			31058: outdata = 32'd34478;
			31059: outdata = 32'd34477;
			31060: outdata = 32'd34476;
			31061: outdata = 32'd34475;
			31062: outdata = 32'd34474;
			31063: outdata = 32'd34473;
			31064: outdata = 32'd34472;
			31065: outdata = 32'd34471;
			31066: outdata = 32'd34470;
			31067: outdata = 32'd34469;
			31068: outdata = 32'd34468;
			31069: outdata = 32'd34467;
			31070: outdata = 32'd34466;
			31071: outdata = 32'd34465;
			31072: outdata = 32'd34464;
			31073: outdata = 32'd34463;
			31074: outdata = 32'd34462;
			31075: outdata = 32'd34461;
			31076: outdata = 32'd34460;
			31077: outdata = 32'd34459;
			31078: outdata = 32'd34458;
			31079: outdata = 32'd34457;
			31080: outdata = 32'd34456;
			31081: outdata = 32'd34455;
			31082: outdata = 32'd34454;
			31083: outdata = 32'd34453;
			31084: outdata = 32'd34452;
			31085: outdata = 32'd34451;
			31086: outdata = 32'd34450;
			31087: outdata = 32'd34449;
			31088: outdata = 32'd34448;
			31089: outdata = 32'd34447;
			31090: outdata = 32'd34446;
			31091: outdata = 32'd34445;
			31092: outdata = 32'd34444;
			31093: outdata = 32'd34443;
			31094: outdata = 32'd34442;
			31095: outdata = 32'd34441;
			31096: outdata = 32'd34440;
			31097: outdata = 32'd34439;
			31098: outdata = 32'd34438;
			31099: outdata = 32'd34437;
			31100: outdata = 32'd34436;
			31101: outdata = 32'd34435;
			31102: outdata = 32'd34434;
			31103: outdata = 32'd34433;
			31104: outdata = 32'd34432;
			31105: outdata = 32'd34431;
			31106: outdata = 32'd34430;
			31107: outdata = 32'd34429;
			31108: outdata = 32'd34428;
			31109: outdata = 32'd34427;
			31110: outdata = 32'd34426;
			31111: outdata = 32'd34425;
			31112: outdata = 32'd34424;
			31113: outdata = 32'd34423;
			31114: outdata = 32'd34422;
			31115: outdata = 32'd34421;
			31116: outdata = 32'd34420;
			31117: outdata = 32'd34419;
			31118: outdata = 32'd34418;
			31119: outdata = 32'd34417;
			31120: outdata = 32'd34416;
			31121: outdata = 32'd34415;
			31122: outdata = 32'd34414;
			31123: outdata = 32'd34413;
			31124: outdata = 32'd34412;
			31125: outdata = 32'd34411;
			31126: outdata = 32'd34410;
			31127: outdata = 32'd34409;
			31128: outdata = 32'd34408;
			31129: outdata = 32'd34407;
			31130: outdata = 32'd34406;
			31131: outdata = 32'd34405;
			31132: outdata = 32'd34404;
			31133: outdata = 32'd34403;
			31134: outdata = 32'd34402;
			31135: outdata = 32'd34401;
			31136: outdata = 32'd34400;
			31137: outdata = 32'd34399;
			31138: outdata = 32'd34398;
			31139: outdata = 32'd34397;
			31140: outdata = 32'd34396;
			31141: outdata = 32'd34395;
			31142: outdata = 32'd34394;
			31143: outdata = 32'd34393;
			31144: outdata = 32'd34392;
			31145: outdata = 32'd34391;
			31146: outdata = 32'd34390;
			31147: outdata = 32'd34389;
			31148: outdata = 32'd34388;
			31149: outdata = 32'd34387;
			31150: outdata = 32'd34386;
			31151: outdata = 32'd34385;
			31152: outdata = 32'd34384;
			31153: outdata = 32'd34383;
			31154: outdata = 32'd34382;
			31155: outdata = 32'd34381;
			31156: outdata = 32'd34380;
			31157: outdata = 32'd34379;
			31158: outdata = 32'd34378;
			31159: outdata = 32'd34377;
			31160: outdata = 32'd34376;
			31161: outdata = 32'd34375;
			31162: outdata = 32'd34374;
			31163: outdata = 32'd34373;
			31164: outdata = 32'd34372;
			31165: outdata = 32'd34371;
			31166: outdata = 32'd34370;
			31167: outdata = 32'd34369;
			31168: outdata = 32'd34368;
			31169: outdata = 32'd34367;
			31170: outdata = 32'd34366;
			31171: outdata = 32'd34365;
			31172: outdata = 32'd34364;
			31173: outdata = 32'd34363;
			31174: outdata = 32'd34362;
			31175: outdata = 32'd34361;
			31176: outdata = 32'd34360;
			31177: outdata = 32'd34359;
			31178: outdata = 32'd34358;
			31179: outdata = 32'd34357;
			31180: outdata = 32'd34356;
			31181: outdata = 32'd34355;
			31182: outdata = 32'd34354;
			31183: outdata = 32'd34353;
			31184: outdata = 32'd34352;
			31185: outdata = 32'd34351;
			31186: outdata = 32'd34350;
			31187: outdata = 32'd34349;
			31188: outdata = 32'd34348;
			31189: outdata = 32'd34347;
			31190: outdata = 32'd34346;
			31191: outdata = 32'd34345;
			31192: outdata = 32'd34344;
			31193: outdata = 32'd34343;
			31194: outdata = 32'd34342;
			31195: outdata = 32'd34341;
			31196: outdata = 32'd34340;
			31197: outdata = 32'd34339;
			31198: outdata = 32'd34338;
			31199: outdata = 32'd34337;
			31200: outdata = 32'd34336;
			31201: outdata = 32'd34335;
			31202: outdata = 32'd34334;
			31203: outdata = 32'd34333;
			31204: outdata = 32'd34332;
			31205: outdata = 32'd34331;
			31206: outdata = 32'd34330;
			31207: outdata = 32'd34329;
			31208: outdata = 32'd34328;
			31209: outdata = 32'd34327;
			31210: outdata = 32'd34326;
			31211: outdata = 32'd34325;
			31212: outdata = 32'd34324;
			31213: outdata = 32'd34323;
			31214: outdata = 32'd34322;
			31215: outdata = 32'd34321;
			31216: outdata = 32'd34320;
			31217: outdata = 32'd34319;
			31218: outdata = 32'd34318;
			31219: outdata = 32'd34317;
			31220: outdata = 32'd34316;
			31221: outdata = 32'd34315;
			31222: outdata = 32'd34314;
			31223: outdata = 32'd34313;
			31224: outdata = 32'd34312;
			31225: outdata = 32'd34311;
			31226: outdata = 32'd34310;
			31227: outdata = 32'd34309;
			31228: outdata = 32'd34308;
			31229: outdata = 32'd34307;
			31230: outdata = 32'd34306;
			31231: outdata = 32'd34305;
			31232: outdata = 32'd34304;
			31233: outdata = 32'd34303;
			31234: outdata = 32'd34302;
			31235: outdata = 32'd34301;
			31236: outdata = 32'd34300;
			31237: outdata = 32'd34299;
			31238: outdata = 32'd34298;
			31239: outdata = 32'd34297;
			31240: outdata = 32'd34296;
			31241: outdata = 32'd34295;
			31242: outdata = 32'd34294;
			31243: outdata = 32'd34293;
			31244: outdata = 32'd34292;
			31245: outdata = 32'd34291;
			31246: outdata = 32'd34290;
			31247: outdata = 32'd34289;
			31248: outdata = 32'd34288;
			31249: outdata = 32'd34287;
			31250: outdata = 32'd34286;
			31251: outdata = 32'd34285;
			31252: outdata = 32'd34284;
			31253: outdata = 32'd34283;
			31254: outdata = 32'd34282;
			31255: outdata = 32'd34281;
			31256: outdata = 32'd34280;
			31257: outdata = 32'd34279;
			31258: outdata = 32'd34278;
			31259: outdata = 32'd34277;
			31260: outdata = 32'd34276;
			31261: outdata = 32'd34275;
			31262: outdata = 32'd34274;
			31263: outdata = 32'd34273;
			31264: outdata = 32'd34272;
			31265: outdata = 32'd34271;
			31266: outdata = 32'd34270;
			31267: outdata = 32'd34269;
			31268: outdata = 32'd34268;
			31269: outdata = 32'd34267;
			31270: outdata = 32'd34266;
			31271: outdata = 32'd34265;
			31272: outdata = 32'd34264;
			31273: outdata = 32'd34263;
			31274: outdata = 32'd34262;
			31275: outdata = 32'd34261;
			31276: outdata = 32'd34260;
			31277: outdata = 32'd34259;
			31278: outdata = 32'd34258;
			31279: outdata = 32'd34257;
			31280: outdata = 32'd34256;
			31281: outdata = 32'd34255;
			31282: outdata = 32'd34254;
			31283: outdata = 32'd34253;
			31284: outdata = 32'd34252;
			31285: outdata = 32'd34251;
			31286: outdata = 32'd34250;
			31287: outdata = 32'd34249;
			31288: outdata = 32'd34248;
			31289: outdata = 32'd34247;
			31290: outdata = 32'd34246;
			31291: outdata = 32'd34245;
			31292: outdata = 32'd34244;
			31293: outdata = 32'd34243;
			31294: outdata = 32'd34242;
			31295: outdata = 32'd34241;
			31296: outdata = 32'd34240;
			31297: outdata = 32'd34239;
			31298: outdata = 32'd34238;
			31299: outdata = 32'd34237;
			31300: outdata = 32'd34236;
			31301: outdata = 32'd34235;
			31302: outdata = 32'd34234;
			31303: outdata = 32'd34233;
			31304: outdata = 32'd34232;
			31305: outdata = 32'd34231;
			31306: outdata = 32'd34230;
			31307: outdata = 32'd34229;
			31308: outdata = 32'd34228;
			31309: outdata = 32'd34227;
			31310: outdata = 32'd34226;
			31311: outdata = 32'd34225;
			31312: outdata = 32'd34224;
			31313: outdata = 32'd34223;
			31314: outdata = 32'd34222;
			31315: outdata = 32'd34221;
			31316: outdata = 32'd34220;
			31317: outdata = 32'd34219;
			31318: outdata = 32'd34218;
			31319: outdata = 32'd34217;
			31320: outdata = 32'd34216;
			31321: outdata = 32'd34215;
			31322: outdata = 32'd34214;
			31323: outdata = 32'd34213;
			31324: outdata = 32'd34212;
			31325: outdata = 32'd34211;
			31326: outdata = 32'd34210;
			31327: outdata = 32'd34209;
			31328: outdata = 32'd34208;
			31329: outdata = 32'd34207;
			31330: outdata = 32'd34206;
			31331: outdata = 32'd34205;
			31332: outdata = 32'd34204;
			31333: outdata = 32'd34203;
			31334: outdata = 32'd34202;
			31335: outdata = 32'd34201;
			31336: outdata = 32'd34200;
			31337: outdata = 32'd34199;
			31338: outdata = 32'd34198;
			31339: outdata = 32'd34197;
			31340: outdata = 32'd34196;
			31341: outdata = 32'd34195;
			31342: outdata = 32'd34194;
			31343: outdata = 32'd34193;
			31344: outdata = 32'd34192;
			31345: outdata = 32'd34191;
			31346: outdata = 32'd34190;
			31347: outdata = 32'd34189;
			31348: outdata = 32'd34188;
			31349: outdata = 32'd34187;
			31350: outdata = 32'd34186;
			31351: outdata = 32'd34185;
			31352: outdata = 32'd34184;
			31353: outdata = 32'd34183;
			31354: outdata = 32'd34182;
			31355: outdata = 32'd34181;
			31356: outdata = 32'd34180;
			31357: outdata = 32'd34179;
			31358: outdata = 32'd34178;
			31359: outdata = 32'd34177;
			31360: outdata = 32'd34176;
			31361: outdata = 32'd34175;
			31362: outdata = 32'd34174;
			31363: outdata = 32'd34173;
			31364: outdata = 32'd34172;
			31365: outdata = 32'd34171;
			31366: outdata = 32'd34170;
			31367: outdata = 32'd34169;
			31368: outdata = 32'd34168;
			31369: outdata = 32'd34167;
			31370: outdata = 32'd34166;
			31371: outdata = 32'd34165;
			31372: outdata = 32'd34164;
			31373: outdata = 32'd34163;
			31374: outdata = 32'd34162;
			31375: outdata = 32'd34161;
			31376: outdata = 32'd34160;
			31377: outdata = 32'd34159;
			31378: outdata = 32'd34158;
			31379: outdata = 32'd34157;
			31380: outdata = 32'd34156;
			31381: outdata = 32'd34155;
			31382: outdata = 32'd34154;
			31383: outdata = 32'd34153;
			31384: outdata = 32'd34152;
			31385: outdata = 32'd34151;
			31386: outdata = 32'd34150;
			31387: outdata = 32'd34149;
			31388: outdata = 32'd34148;
			31389: outdata = 32'd34147;
			31390: outdata = 32'd34146;
			31391: outdata = 32'd34145;
			31392: outdata = 32'd34144;
			31393: outdata = 32'd34143;
			31394: outdata = 32'd34142;
			31395: outdata = 32'd34141;
			31396: outdata = 32'd34140;
			31397: outdata = 32'd34139;
			31398: outdata = 32'd34138;
			31399: outdata = 32'd34137;
			31400: outdata = 32'd34136;
			31401: outdata = 32'd34135;
			31402: outdata = 32'd34134;
			31403: outdata = 32'd34133;
			31404: outdata = 32'd34132;
			31405: outdata = 32'd34131;
			31406: outdata = 32'd34130;
			31407: outdata = 32'd34129;
			31408: outdata = 32'd34128;
			31409: outdata = 32'd34127;
			31410: outdata = 32'd34126;
			31411: outdata = 32'd34125;
			31412: outdata = 32'd34124;
			31413: outdata = 32'd34123;
			31414: outdata = 32'd34122;
			31415: outdata = 32'd34121;
			31416: outdata = 32'd34120;
			31417: outdata = 32'd34119;
			31418: outdata = 32'd34118;
			31419: outdata = 32'd34117;
			31420: outdata = 32'd34116;
			31421: outdata = 32'd34115;
			31422: outdata = 32'd34114;
			31423: outdata = 32'd34113;
			31424: outdata = 32'd34112;
			31425: outdata = 32'd34111;
			31426: outdata = 32'd34110;
			31427: outdata = 32'd34109;
			31428: outdata = 32'd34108;
			31429: outdata = 32'd34107;
			31430: outdata = 32'd34106;
			31431: outdata = 32'd34105;
			31432: outdata = 32'd34104;
			31433: outdata = 32'd34103;
			31434: outdata = 32'd34102;
			31435: outdata = 32'd34101;
			31436: outdata = 32'd34100;
			31437: outdata = 32'd34099;
			31438: outdata = 32'd34098;
			31439: outdata = 32'd34097;
			31440: outdata = 32'd34096;
			31441: outdata = 32'd34095;
			31442: outdata = 32'd34094;
			31443: outdata = 32'd34093;
			31444: outdata = 32'd34092;
			31445: outdata = 32'd34091;
			31446: outdata = 32'd34090;
			31447: outdata = 32'd34089;
			31448: outdata = 32'd34088;
			31449: outdata = 32'd34087;
			31450: outdata = 32'd34086;
			31451: outdata = 32'd34085;
			31452: outdata = 32'd34084;
			31453: outdata = 32'd34083;
			31454: outdata = 32'd34082;
			31455: outdata = 32'd34081;
			31456: outdata = 32'd34080;
			31457: outdata = 32'd34079;
			31458: outdata = 32'd34078;
			31459: outdata = 32'd34077;
			31460: outdata = 32'd34076;
			31461: outdata = 32'd34075;
			31462: outdata = 32'd34074;
			31463: outdata = 32'd34073;
			31464: outdata = 32'd34072;
			31465: outdata = 32'd34071;
			31466: outdata = 32'd34070;
			31467: outdata = 32'd34069;
			31468: outdata = 32'd34068;
			31469: outdata = 32'd34067;
			31470: outdata = 32'd34066;
			31471: outdata = 32'd34065;
			31472: outdata = 32'd34064;
			31473: outdata = 32'd34063;
			31474: outdata = 32'd34062;
			31475: outdata = 32'd34061;
			31476: outdata = 32'd34060;
			31477: outdata = 32'd34059;
			31478: outdata = 32'd34058;
			31479: outdata = 32'd34057;
			31480: outdata = 32'd34056;
			31481: outdata = 32'd34055;
			31482: outdata = 32'd34054;
			31483: outdata = 32'd34053;
			31484: outdata = 32'd34052;
			31485: outdata = 32'd34051;
			31486: outdata = 32'd34050;
			31487: outdata = 32'd34049;
			31488: outdata = 32'd34048;
			31489: outdata = 32'd34047;
			31490: outdata = 32'd34046;
			31491: outdata = 32'd34045;
			31492: outdata = 32'd34044;
			31493: outdata = 32'd34043;
			31494: outdata = 32'd34042;
			31495: outdata = 32'd34041;
			31496: outdata = 32'd34040;
			31497: outdata = 32'd34039;
			31498: outdata = 32'd34038;
			31499: outdata = 32'd34037;
			31500: outdata = 32'd34036;
			31501: outdata = 32'd34035;
			31502: outdata = 32'd34034;
			31503: outdata = 32'd34033;
			31504: outdata = 32'd34032;
			31505: outdata = 32'd34031;
			31506: outdata = 32'd34030;
			31507: outdata = 32'd34029;
			31508: outdata = 32'd34028;
			31509: outdata = 32'd34027;
			31510: outdata = 32'd34026;
			31511: outdata = 32'd34025;
			31512: outdata = 32'd34024;
			31513: outdata = 32'd34023;
			31514: outdata = 32'd34022;
			31515: outdata = 32'd34021;
			31516: outdata = 32'd34020;
			31517: outdata = 32'd34019;
			31518: outdata = 32'd34018;
			31519: outdata = 32'd34017;
			31520: outdata = 32'd34016;
			31521: outdata = 32'd34015;
			31522: outdata = 32'd34014;
			31523: outdata = 32'd34013;
			31524: outdata = 32'd34012;
			31525: outdata = 32'd34011;
			31526: outdata = 32'd34010;
			31527: outdata = 32'd34009;
			31528: outdata = 32'd34008;
			31529: outdata = 32'd34007;
			31530: outdata = 32'd34006;
			31531: outdata = 32'd34005;
			31532: outdata = 32'd34004;
			31533: outdata = 32'd34003;
			31534: outdata = 32'd34002;
			31535: outdata = 32'd34001;
			31536: outdata = 32'd34000;
			31537: outdata = 32'd33999;
			31538: outdata = 32'd33998;
			31539: outdata = 32'd33997;
			31540: outdata = 32'd33996;
			31541: outdata = 32'd33995;
			31542: outdata = 32'd33994;
			31543: outdata = 32'd33993;
			31544: outdata = 32'd33992;
			31545: outdata = 32'd33991;
			31546: outdata = 32'd33990;
			31547: outdata = 32'd33989;
			31548: outdata = 32'd33988;
			31549: outdata = 32'd33987;
			31550: outdata = 32'd33986;
			31551: outdata = 32'd33985;
			31552: outdata = 32'd33984;
			31553: outdata = 32'd33983;
			31554: outdata = 32'd33982;
			31555: outdata = 32'd33981;
			31556: outdata = 32'd33980;
			31557: outdata = 32'd33979;
			31558: outdata = 32'd33978;
			31559: outdata = 32'd33977;
			31560: outdata = 32'd33976;
			31561: outdata = 32'd33975;
			31562: outdata = 32'd33974;
			31563: outdata = 32'd33973;
			31564: outdata = 32'd33972;
			31565: outdata = 32'd33971;
			31566: outdata = 32'd33970;
			31567: outdata = 32'd33969;
			31568: outdata = 32'd33968;
			31569: outdata = 32'd33967;
			31570: outdata = 32'd33966;
			31571: outdata = 32'd33965;
			31572: outdata = 32'd33964;
			31573: outdata = 32'd33963;
			31574: outdata = 32'd33962;
			31575: outdata = 32'd33961;
			31576: outdata = 32'd33960;
			31577: outdata = 32'd33959;
			31578: outdata = 32'd33958;
			31579: outdata = 32'd33957;
			31580: outdata = 32'd33956;
			31581: outdata = 32'd33955;
			31582: outdata = 32'd33954;
			31583: outdata = 32'd33953;
			31584: outdata = 32'd33952;
			31585: outdata = 32'd33951;
			31586: outdata = 32'd33950;
			31587: outdata = 32'd33949;
			31588: outdata = 32'd33948;
			31589: outdata = 32'd33947;
			31590: outdata = 32'd33946;
			31591: outdata = 32'd33945;
			31592: outdata = 32'd33944;
			31593: outdata = 32'd33943;
			31594: outdata = 32'd33942;
			31595: outdata = 32'd33941;
			31596: outdata = 32'd33940;
			31597: outdata = 32'd33939;
			31598: outdata = 32'd33938;
			31599: outdata = 32'd33937;
			31600: outdata = 32'd33936;
			31601: outdata = 32'd33935;
			31602: outdata = 32'd33934;
			31603: outdata = 32'd33933;
			31604: outdata = 32'd33932;
			31605: outdata = 32'd33931;
			31606: outdata = 32'd33930;
			31607: outdata = 32'd33929;
			31608: outdata = 32'd33928;
			31609: outdata = 32'd33927;
			31610: outdata = 32'd33926;
			31611: outdata = 32'd33925;
			31612: outdata = 32'd33924;
			31613: outdata = 32'd33923;
			31614: outdata = 32'd33922;
			31615: outdata = 32'd33921;
			31616: outdata = 32'd33920;
			31617: outdata = 32'd33919;
			31618: outdata = 32'd33918;
			31619: outdata = 32'd33917;
			31620: outdata = 32'd33916;
			31621: outdata = 32'd33915;
			31622: outdata = 32'd33914;
			31623: outdata = 32'd33913;
			31624: outdata = 32'd33912;
			31625: outdata = 32'd33911;
			31626: outdata = 32'd33910;
			31627: outdata = 32'd33909;
			31628: outdata = 32'd33908;
			31629: outdata = 32'd33907;
			31630: outdata = 32'd33906;
			31631: outdata = 32'd33905;
			31632: outdata = 32'd33904;
			31633: outdata = 32'd33903;
			31634: outdata = 32'd33902;
			31635: outdata = 32'd33901;
			31636: outdata = 32'd33900;
			31637: outdata = 32'd33899;
			31638: outdata = 32'd33898;
			31639: outdata = 32'd33897;
			31640: outdata = 32'd33896;
			31641: outdata = 32'd33895;
			31642: outdata = 32'd33894;
			31643: outdata = 32'd33893;
			31644: outdata = 32'd33892;
			31645: outdata = 32'd33891;
			31646: outdata = 32'd33890;
			31647: outdata = 32'd33889;
			31648: outdata = 32'd33888;
			31649: outdata = 32'd33887;
			31650: outdata = 32'd33886;
			31651: outdata = 32'd33885;
			31652: outdata = 32'd33884;
			31653: outdata = 32'd33883;
			31654: outdata = 32'd33882;
			31655: outdata = 32'd33881;
			31656: outdata = 32'd33880;
			31657: outdata = 32'd33879;
			31658: outdata = 32'd33878;
			31659: outdata = 32'd33877;
			31660: outdata = 32'd33876;
			31661: outdata = 32'd33875;
			31662: outdata = 32'd33874;
			31663: outdata = 32'd33873;
			31664: outdata = 32'd33872;
			31665: outdata = 32'd33871;
			31666: outdata = 32'd33870;
			31667: outdata = 32'd33869;
			31668: outdata = 32'd33868;
			31669: outdata = 32'd33867;
			31670: outdata = 32'd33866;
			31671: outdata = 32'd33865;
			31672: outdata = 32'd33864;
			31673: outdata = 32'd33863;
			31674: outdata = 32'd33862;
			31675: outdata = 32'd33861;
			31676: outdata = 32'd33860;
			31677: outdata = 32'd33859;
			31678: outdata = 32'd33858;
			31679: outdata = 32'd33857;
			31680: outdata = 32'd33856;
			31681: outdata = 32'd33855;
			31682: outdata = 32'd33854;
			31683: outdata = 32'd33853;
			31684: outdata = 32'd33852;
			31685: outdata = 32'd33851;
			31686: outdata = 32'd33850;
			31687: outdata = 32'd33849;
			31688: outdata = 32'd33848;
			31689: outdata = 32'd33847;
			31690: outdata = 32'd33846;
			31691: outdata = 32'd33845;
			31692: outdata = 32'd33844;
			31693: outdata = 32'd33843;
			31694: outdata = 32'd33842;
			31695: outdata = 32'd33841;
			31696: outdata = 32'd33840;
			31697: outdata = 32'd33839;
			31698: outdata = 32'd33838;
			31699: outdata = 32'd33837;
			31700: outdata = 32'd33836;
			31701: outdata = 32'd33835;
			31702: outdata = 32'd33834;
			31703: outdata = 32'd33833;
			31704: outdata = 32'd33832;
			31705: outdata = 32'd33831;
			31706: outdata = 32'd33830;
			31707: outdata = 32'd33829;
			31708: outdata = 32'd33828;
			31709: outdata = 32'd33827;
			31710: outdata = 32'd33826;
			31711: outdata = 32'd33825;
			31712: outdata = 32'd33824;
			31713: outdata = 32'd33823;
			31714: outdata = 32'd33822;
			31715: outdata = 32'd33821;
			31716: outdata = 32'd33820;
			31717: outdata = 32'd33819;
			31718: outdata = 32'd33818;
			31719: outdata = 32'd33817;
			31720: outdata = 32'd33816;
			31721: outdata = 32'd33815;
			31722: outdata = 32'd33814;
			31723: outdata = 32'd33813;
			31724: outdata = 32'd33812;
			31725: outdata = 32'd33811;
			31726: outdata = 32'd33810;
			31727: outdata = 32'd33809;
			31728: outdata = 32'd33808;
			31729: outdata = 32'd33807;
			31730: outdata = 32'd33806;
			31731: outdata = 32'd33805;
			31732: outdata = 32'd33804;
			31733: outdata = 32'd33803;
			31734: outdata = 32'd33802;
			31735: outdata = 32'd33801;
			31736: outdata = 32'd33800;
			31737: outdata = 32'd33799;
			31738: outdata = 32'd33798;
			31739: outdata = 32'd33797;
			31740: outdata = 32'd33796;
			31741: outdata = 32'd33795;
			31742: outdata = 32'd33794;
			31743: outdata = 32'd33793;
			31744: outdata = 32'd33792;
			31745: outdata = 32'd33791;
			31746: outdata = 32'd33790;
			31747: outdata = 32'd33789;
			31748: outdata = 32'd33788;
			31749: outdata = 32'd33787;
			31750: outdata = 32'd33786;
			31751: outdata = 32'd33785;
			31752: outdata = 32'd33784;
			31753: outdata = 32'd33783;
			31754: outdata = 32'd33782;
			31755: outdata = 32'd33781;
			31756: outdata = 32'd33780;
			31757: outdata = 32'd33779;
			31758: outdata = 32'd33778;
			31759: outdata = 32'd33777;
			31760: outdata = 32'd33776;
			31761: outdata = 32'd33775;
			31762: outdata = 32'd33774;
			31763: outdata = 32'd33773;
			31764: outdata = 32'd33772;
			31765: outdata = 32'd33771;
			31766: outdata = 32'd33770;
			31767: outdata = 32'd33769;
			31768: outdata = 32'd33768;
			31769: outdata = 32'd33767;
			31770: outdata = 32'd33766;
			31771: outdata = 32'd33765;
			31772: outdata = 32'd33764;
			31773: outdata = 32'd33763;
			31774: outdata = 32'd33762;
			31775: outdata = 32'd33761;
			31776: outdata = 32'd33760;
			31777: outdata = 32'd33759;
			31778: outdata = 32'd33758;
			31779: outdata = 32'd33757;
			31780: outdata = 32'd33756;
			31781: outdata = 32'd33755;
			31782: outdata = 32'd33754;
			31783: outdata = 32'd33753;
			31784: outdata = 32'd33752;
			31785: outdata = 32'd33751;
			31786: outdata = 32'd33750;
			31787: outdata = 32'd33749;
			31788: outdata = 32'd33748;
			31789: outdata = 32'd33747;
			31790: outdata = 32'd33746;
			31791: outdata = 32'd33745;
			31792: outdata = 32'd33744;
			31793: outdata = 32'd33743;
			31794: outdata = 32'd33742;
			31795: outdata = 32'd33741;
			31796: outdata = 32'd33740;
			31797: outdata = 32'd33739;
			31798: outdata = 32'd33738;
			31799: outdata = 32'd33737;
			31800: outdata = 32'd33736;
			31801: outdata = 32'd33735;
			31802: outdata = 32'd33734;
			31803: outdata = 32'd33733;
			31804: outdata = 32'd33732;
			31805: outdata = 32'd33731;
			31806: outdata = 32'd33730;
			31807: outdata = 32'd33729;
			31808: outdata = 32'd33728;
			31809: outdata = 32'd33727;
			31810: outdata = 32'd33726;
			31811: outdata = 32'd33725;
			31812: outdata = 32'd33724;
			31813: outdata = 32'd33723;
			31814: outdata = 32'd33722;
			31815: outdata = 32'd33721;
			31816: outdata = 32'd33720;
			31817: outdata = 32'd33719;
			31818: outdata = 32'd33718;
			31819: outdata = 32'd33717;
			31820: outdata = 32'd33716;
			31821: outdata = 32'd33715;
			31822: outdata = 32'd33714;
			31823: outdata = 32'd33713;
			31824: outdata = 32'd33712;
			31825: outdata = 32'd33711;
			31826: outdata = 32'd33710;
			31827: outdata = 32'd33709;
			31828: outdata = 32'd33708;
			31829: outdata = 32'd33707;
			31830: outdata = 32'd33706;
			31831: outdata = 32'd33705;
			31832: outdata = 32'd33704;
			31833: outdata = 32'd33703;
			31834: outdata = 32'd33702;
			31835: outdata = 32'd33701;
			31836: outdata = 32'd33700;
			31837: outdata = 32'd33699;
			31838: outdata = 32'd33698;
			31839: outdata = 32'd33697;
			31840: outdata = 32'd33696;
			31841: outdata = 32'd33695;
			31842: outdata = 32'd33694;
			31843: outdata = 32'd33693;
			31844: outdata = 32'd33692;
			31845: outdata = 32'd33691;
			31846: outdata = 32'd33690;
			31847: outdata = 32'd33689;
			31848: outdata = 32'd33688;
			31849: outdata = 32'd33687;
			31850: outdata = 32'd33686;
			31851: outdata = 32'd33685;
			31852: outdata = 32'd33684;
			31853: outdata = 32'd33683;
			31854: outdata = 32'd33682;
			31855: outdata = 32'd33681;
			31856: outdata = 32'd33680;
			31857: outdata = 32'd33679;
			31858: outdata = 32'd33678;
			31859: outdata = 32'd33677;
			31860: outdata = 32'd33676;
			31861: outdata = 32'd33675;
			31862: outdata = 32'd33674;
			31863: outdata = 32'd33673;
			31864: outdata = 32'd33672;
			31865: outdata = 32'd33671;
			31866: outdata = 32'd33670;
			31867: outdata = 32'd33669;
			31868: outdata = 32'd33668;
			31869: outdata = 32'd33667;
			31870: outdata = 32'd33666;
			31871: outdata = 32'd33665;
			31872: outdata = 32'd33664;
			31873: outdata = 32'd33663;
			31874: outdata = 32'd33662;
			31875: outdata = 32'd33661;
			31876: outdata = 32'd33660;
			31877: outdata = 32'd33659;
			31878: outdata = 32'd33658;
			31879: outdata = 32'd33657;
			31880: outdata = 32'd33656;
			31881: outdata = 32'd33655;
			31882: outdata = 32'd33654;
			31883: outdata = 32'd33653;
			31884: outdata = 32'd33652;
			31885: outdata = 32'd33651;
			31886: outdata = 32'd33650;
			31887: outdata = 32'd33649;
			31888: outdata = 32'd33648;
			31889: outdata = 32'd33647;
			31890: outdata = 32'd33646;
			31891: outdata = 32'd33645;
			31892: outdata = 32'd33644;
			31893: outdata = 32'd33643;
			31894: outdata = 32'd33642;
			31895: outdata = 32'd33641;
			31896: outdata = 32'd33640;
			31897: outdata = 32'd33639;
			31898: outdata = 32'd33638;
			31899: outdata = 32'd33637;
			31900: outdata = 32'd33636;
			31901: outdata = 32'd33635;
			31902: outdata = 32'd33634;
			31903: outdata = 32'd33633;
			31904: outdata = 32'd33632;
			31905: outdata = 32'd33631;
			31906: outdata = 32'd33630;
			31907: outdata = 32'd33629;
			31908: outdata = 32'd33628;
			31909: outdata = 32'd33627;
			31910: outdata = 32'd33626;
			31911: outdata = 32'd33625;
			31912: outdata = 32'd33624;
			31913: outdata = 32'd33623;
			31914: outdata = 32'd33622;
			31915: outdata = 32'd33621;
			31916: outdata = 32'd33620;
			31917: outdata = 32'd33619;
			31918: outdata = 32'd33618;
			31919: outdata = 32'd33617;
			31920: outdata = 32'd33616;
			31921: outdata = 32'd33615;
			31922: outdata = 32'd33614;
			31923: outdata = 32'd33613;
			31924: outdata = 32'd33612;
			31925: outdata = 32'd33611;
			31926: outdata = 32'd33610;
			31927: outdata = 32'd33609;
			31928: outdata = 32'd33608;
			31929: outdata = 32'd33607;
			31930: outdata = 32'd33606;
			31931: outdata = 32'd33605;
			31932: outdata = 32'd33604;
			31933: outdata = 32'd33603;
			31934: outdata = 32'd33602;
			31935: outdata = 32'd33601;
			31936: outdata = 32'd33600;
			31937: outdata = 32'd33599;
			31938: outdata = 32'd33598;
			31939: outdata = 32'd33597;
			31940: outdata = 32'd33596;
			31941: outdata = 32'd33595;
			31942: outdata = 32'd33594;
			31943: outdata = 32'd33593;
			31944: outdata = 32'd33592;
			31945: outdata = 32'd33591;
			31946: outdata = 32'd33590;
			31947: outdata = 32'd33589;
			31948: outdata = 32'd33588;
			31949: outdata = 32'd33587;
			31950: outdata = 32'd33586;
			31951: outdata = 32'd33585;
			31952: outdata = 32'd33584;
			31953: outdata = 32'd33583;
			31954: outdata = 32'd33582;
			31955: outdata = 32'd33581;
			31956: outdata = 32'd33580;
			31957: outdata = 32'd33579;
			31958: outdata = 32'd33578;
			31959: outdata = 32'd33577;
			31960: outdata = 32'd33576;
			31961: outdata = 32'd33575;
			31962: outdata = 32'd33574;
			31963: outdata = 32'd33573;
			31964: outdata = 32'd33572;
			31965: outdata = 32'd33571;
			31966: outdata = 32'd33570;
			31967: outdata = 32'd33569;
			31968: outdata = 32'd33568;
			31969: outdata = 32'd33567;
			31970: outdata = 32'd33566;
			31971: outdata = 32'd33565;
			31972: outdata = 32'd33564;
			31973: outdata = 32'd33563;
			31974: outdata = 32'd33562;
			31975: outdata = 32'd33561;
			31976: outdata = 32'd33560;
			31977: outdata = 32'd33559;
			31978: outdata = 32'd33558;
			31979: outdata = 32'd33557;
			31980: outdata = 32'd33556;
			31981: outdata = 32'd33555;
			31982: outdata = 32'd33554;
			31983: outdata = 32'd33553;
			31984: outdata = 32'd33552;
			31985: outdata = 32'd33551;
			31986: outdata = 32'd33550;
			31987: outdata = 32'd33549;
			31988: outdata = 32'd33548;
			31989: outdata = 32'd33547;
			31990: outdata = 32'd33546;
			31991: outdata = 32'd33545;
			31992: outdata = 32'd33544;
			31993: outdata = 32'd33543;
			31994: outdata = 32'd33542;
			31995: outdata = 32'd33541;
			31996: outdata = 32'd33540;
			31997: outdata = 32'd33539;
			31998: outdata = 32'd33538;
			31999: outdata = 32'd33537;
			32000: outdata = 32'd33536;
			32001: outdata = 32'd33535;
			32002: outdata = 32'd33534;
			32003: outdata = 32'd33533;
			32004: outdata = 32'd33532;
			32005: outdata = 32'd33531;
			32006: outdata = 32'd33530;
			32007: outdata = 32'd33529;
			32008: outdata = 32'd33528;
			32009: outdata = 32'd33527;
			32010: outdata = 32'd33526;
			32011: outdata = 32'd33525;
			32012: outdata = 32'd33524;
			32013: outdata = 32'd33523;
			32014: outdata = 32'd33522;
			32015: outdata = 32'd33521;
			32016: outdata = 32'd33520;
			32017: outdata = 32'd33519;
			32018: outdata = 32'd33518;
			32019: outdata = 32'd33517;
			32020: outdata = 32'd33516;
			32021: outdata = 32'd33515;
			32022: outdata = 32'd33514;
			32023: outdata = 32'd33513;
			32024: outdata = 32'd33512;
			32025: outdata = 32'd33511;
			32026: outdata = 32'd33510;
			32027: outdata = 32'd33509;
			32028: outdata = 32'd33508;
			32029: outdata = 32'd33507;
			32030: outdata = 32'd33506;
			32031: outdata = 32'd33505;
			32032: outdata = 32'd33504;
			32033: outdata = 32'd33503;
			32034: outdata = 32'd33502;
			32035: outdata = 32'd33501;
			32036: outdata = 32'd33500;
			32037: outdata = 32'd33499;
			32038: outdata = 32'd33498;
			32039: outdata = 32'd33497;
			32040: outdata = 32'd33496;
			32041: outdata = 32'd33495;
			32042: outdata = 32'd33494;
			32043: outdata = 32'd33493;
			32044: outdata = 32'd33492;
			32045: outdata = 32'd33491;
			32046: outdata = 32'd33490;
			32047: outdata = 32'd33489;
			32048: outdata = 32'd33488;
			32049: outdata = 32'd33487;
			32050: outdata = 32'd33486;
			32051: outdata = 32'd33485;
			32052: outdata = 32'd33484;
			32053: outdata = 32'd33483;
			32054: outdata = 32'd33482;
			32055: outdata = 32'd33481;
			32056: outdata = 32'd33480;
			32057: outdata = 32'd33479;
			32058: outdata = 32'd33478;
			32059: outdata = 32'd33477;
			32060: outdata = 32'd33476;
			32061: outdata = 32'd33475;
			32062: outdata = 32'd33474;
			32063: outdata = 32'd33473;
			32064: outdata = 32'd33472;
			32065: outdata = 32'd33471;
			32066: outdata = 32'd33470;
			32067: outdata = 32'd33469;
			32068: outdata = 32'd33468;
			32069: outdata = 32'd33467;
			32070: outdata = 32'd33466;
			32071: outdata = 32'd33465;
			32072: outdata = 32'd33464;
			32073: outdata = 32'd33463;
			32074: outdata = 32'd33462;
			32075: outdata = 32'd33461;
			32076: outdata = 32'd33460;
			32077: outdata = 32'd33459;
			32078: outdata = 32'd33458;
			32079: outdata = 32'd33457;
			32080: outdata = 32'd33456;
			32081: outdata = 32'd33455;
			32082: outdata = 32'd33454;
			32083: outdata = 32'd33453;
			32084: outdata = 32'd33452;
			32085: outdata = 32'd33451;
			32086: outdata = 32'd33450;
			32087: outdata = 32'd33449;
			32088: outdata = 32'd33448;
			32089: outdata = 32'd33447;
			32090: outdata = 32'd33446;
			32091: outdata = 32'd33445;
			32092: outdata = 32'd33444;
			32093: outdata = 32'd33443;
			32094: outdata = 32'd33442;
			32095: outdata = 32'd33441;
			32096: outdata = 32'd33440;
			32097: outdata = 32'd33439;
			32098: outdata = 32'd33438;
			32099: outdata = 32'd33437;
			32100: outdata = 32'd33436;
			32101: outdata = 32'd33435;
			32102: outdata = 32'd33434;
			32103: outdata = 32'd33433;
			32104: outdata = 32'd33432;
			32105: outdata = 32'd33431;
			32106: outdata = 32'd33430;
			32107: outdata = 32'd33429;
			32108: outdata = 32'd33428;
			32109: outdata = 32'd33427;
			32110: outdata = 32'd33426;
			32111: outdata = 32'd33425;
			32112: outdata = 32'd33424;
			32113: outdata = 32'd33423;
			32114: outdata = 32'd33422;
			32115: outdata = 32'd33421;
			32116: outdata = 32'd33420;
			32117: outdata = 32'd33419;
			32118: outdata = 32'd33418;
			32119: outdata = 32'd33417;
			32120: outdata = 32'd33416;
			32121: outdata = 32'd33415;
			32122: outdata = 32'd33414;
			32123: outdata = 32'd33413;
			32124: outdata = 32'd33412;
			32125: outdata = 32'd33411;
			32126: outdata = 32'd33410;
			32127: outdata = 32'd33409;
			32128: outdata = 32'd33408;
			32129: outdata = 32'd33407;
			32130: outdata = 32'd33406;
			32131: outdata = 32'd33405;
			32132: outdata = 32'd33404;
			32133: outdata = 32'd33403;
			32134: outdata = 32'd33402;
			32135: outdata = 32'd33401;
			32136: outdata = 32'd33400;
			32137: outdata = 32'd33399;
			32138: outdata = 32'd33398;
			32139: outdata = 32'd33397;
			32140: outdata = 32'd33396;
			32141: outdata = 32'd33395;
			32142: outdata = 32'd33394;
			32143: outdata = 32'd33393;
			32144: outdata = 32'd33392;
			32145: outdata = 32'd33391;
			32146: outdata = 32'd33390;
			32147: outdata = 32'd33389;
			32148: outdata = 32'd33388;
			32149: outdata = 32'd33387;
			32150: outdata = 32'd33386;
			32151: outdata = 32'd33385;
			32152: outdata = 32'd33384;
			32153: outdata = 32'd33383;
			32154: outdata = 32'd33382;
			32155: outdata = 32'd33381;
			32156: outdata = 32'd33380;
			32157: outdata = 32'd33379;
			32158: outdata = 32'd33378;
			32159: outdata = 32'd33377;
			32160: outdata = 32'd33376;
			32161: outdata = 32'd33375;
			32162: outdata = 32'd33374;
			32163: outdata = 32'd33373;
			32164: outdata = 32'd33372;
			32165: outdata = 32'd33371;
			32166: outdata = 32'd33370;
			32167: outdata = 32'd33369;
			32168: outdata = 32'd33368;
			32169: outdata = 32'd33367;
			32170: outdata = 32'd33366;
			32171: outdata = 32'd33365;
			32172: outdata = 32'd33364;
			32173: outdata = 32'd33363;
			32174: outdata = 32'd33362;
			32175: outdata = 32'd33361;
			32176: outdata = 32'd33360;
			32177: outdata = 32'd33359;
			32178: outdata = 32'd33358;
			32179: outdata = 32'd33357;
			32180: outdata = 32'd33356;
			32181: outdata = 32'd33355;
			32182: outdata = 32'd33354;
			32183: outdata = 32'd33353;
			32184: outdata = 32'd33352;
			32185: outdata = 32'd33351;
			32186: outdata = 32'd33350;
			32187: outdata = 32'd33349;
			32188: outdata = 32'd33348;
			32189: outdata = 32'd33347;
			32190: outdata = 32'd33346;
			32191: outdata = 32'd33345;
			32192: outdata = 32'd33344;
			32193: outdata = 32'd33343;
			32194: outdata = 32'd33342;
			32195: outdata = 32'd33341;
			32196: outdata = 32'd33340;
			32197: outdata = 32'd33339;
			32198: outdata = 32'd33338;
			32199: outdata = 32'd33337;
			32200: outdata = 32'd33336;
			32201: outdata = 32'd33335;
			32202: outdata = 32'd33334;
			32203: outdata = 32'd33333;
			32204: outdata = 32'd33332;
			32205: outdata = 32'd33331;
			32206: outdata = 32'd33330;
			32207: outdata = 32'd33329;
			32208: outdata = 32'd33328;
			32209: outdata = 32'd33327;
			32210: outdata = 32'd33326;
			32211: outdata = 32'd33325;
			32212: outdata = 32'd33324;
			32213: outdata = 32'd33323;
			32214: outdata = 32'd33322;
			32215: outdata = 32'd33321;
			32216: outdata = 32'd33320;
			32217: outdata = 32'd33319;
			32218: outdata = 32'd33318;
			32219: outdata = 32'd33317;
			32220: outdata = 32'd33316;
			32221: outdata = 32'd33315;
			32222: outdata = 32'd33314;
			32223: outdata = 32'd33313;
			32224: outdata = 32'd33312;
			32225: outdata = 32'd33311;
			32226: outdata = 32'd33310;
			32227: outdata = 32'd33309;
			32228: outdata = 32'd33308;
			32229: outdata = 32'd33307;
			32230: outdata = 32'd33306;
			32231: outdata = 32'd33305;
			32232: outdata = 32'd33304;
			32233: outdata = 32'd33303;
			32234: outdata = 32'd33302;
			32235: outdata = 32'd33301;
			32236: outdata = 32'd33300;
			32237: outdata = 32'd33299;
			32238: outdata = 32'd33298;
			32239: outdata = 32'd33297;
			32240: outdata = 32'd33296;
			32241: outdata = 32'd33295;
			32242: outdata = 32'd33294;
			32243: outdata = 32'd33293;
			32244: outdata = 32'd33292;
			32245: outdata = 32'd33291;
			32246: outdata = 32'd33290;
			32247: outdata = 32'd33289;
			32248: outdata = 32'd33288;
			32249: outdata = 32'd33287;
			32250: outdata = 32'd33286;
			32251: outdata = 32'd33285;
			32252: outdata = 32'd33284;
			32253: outdata = 32'd33283;
			32254: outdata = 32'd33282;
			32255: outdata = 32'd33281;
			32256: outdata = 32'd33280;
			32257: outdata = 32'd33279;
			32258: outdata = 32'd33278;
			32259: outdata = 32'd33277;
			32260: outdata = 32'd33276;
			32261: outdata = 32'd33275;
			32262: outdata = 32'd33274;
			32263: outdata = 32'd33273;
			32264: outdata = 32'd33272;
			32265: outdata = 32'd33271;
			32266: outdata = 32'd33270;
			32267: outdata = 32'd33269;
			32268: outdata = 32'd33268;
			32269: outdata = 32'd33267;
			32270: outdata = 32'd33266;
			32271: outdata = 32'd33265;
			32272: outdata = 32'd33264;
			32273: outdata = 32'd33263;
			32274: outdata = 32'd33262;
			32275: outdata = 32'd33261;
			32276: outdata = 32'd33260;
			32277: outdata = 32'd33259;
			32278: outdata = 32'd33258;
			32279: outdata = 32'd33257;
			32280: outdata = 32'd33256;
			32281: outdata = 32'd33255;
			32282: outdata = 32'd33254;
			32283: outdata = 32'd33253;
			32284: outdata = 32'd33252;
			32285: outdata = 32'd33251;
			32286: outdata = 32'd33250;
			32287: outdata = 32'd33249;
			32288: outdata = 32'd33248;
			32289: outdata = 32'd33247;
			32290: outdata = 32'd33246;
			32291: outdata = 32'd33245;
			32292: outdata = 32'd33244;
			32293: outdata = 32'd33243;
			32294: outdata = 32'd33242;
			32295: outdata = 32'd33241;
			32296: outdata = 32'd33240;
			32297: outdata = 32'd33239;
			32298: outdata = 32'd33238;
			32299: outdata = 32'd33237;
			32300: outdata = 32'd33236;
			32301: outdata = 32'd33235;
			32302: outdata = 32'd33234;
			32303: outdata = 32'd33233;
			32304: outdata = 32'd33232;
			32305: outdata = 32'd33231;
			32306: outdata = 32'd33230;
			32307: outdata = 32'd33229;
			32308: outdata = 32'd33228;
			32309: outdata = 32'd33227;
			32310: outdata = 32'd33226;
			32311: outdata = 32'd33225;
			32312: outdata = 32'd33224;
			32313: outdata = 32'd33223;
			32314: outdata = 32'd33222;
			32315: outdata = 32'd33221;
			32316: outdata = 32'd33220;
			32317: outdata = 32'd33219;
			32318: outdata = 32'd33218;
			32319: outdata = 32'd33217;
			32320: outdata = 32'd33216;
			32321: outdata = 32'd33215;
			32322: outdata = 32'd33214;
			32323: outdata = 32'd33213;
			32324: outdata = 32'd33212;
			32325: outdata = 32'd33211;
			32326: outdata = 32'd33210;
			32327: outdata = 32'd33209;
			32328: outdata = 32'd33208;
			32329: outdata = 32'd33207;
			32330: outdata = 32'd33206;
			32331: outdata = 32'd33205;
			32332: outdata = 32'd33204;
			32333: outdata = 32'd33203;
			32334: outdata = 32'd33202;
			32335: outdata = 32'd33201;
			32336: outdata = 32'd33200;
			32337: outdata = 32'd33199;
			32338: outdata = 32'd33198;
			32339: outdata = 32'd33197;
			32340: outdata = 32'd33196;
			32341: outdata = 32'd33195;
			32342: outdata = 32'd33194;
			32343: outdata = 32'd33193;
			32344: outdata = 32'd33192;
			32345: outdata = 32'd33191;
			32346: outdata = 32'd33190;
			32347: outdata = 32'd33189;
			32348: outdata = 32'd33188;
			32349: outdata = 32'd33187;
			32350: outdata = 32'd33186;
			32351: outdata = 32'd33185;
			32352: outdata = 32'd33184;
			32353: outdata = 32'd33183;
			32354: outdata = 32'd33182;
			32355: outdata = 32'd33181;
			32356: outdata = 32'd33180;
			32357: outdata = 32'd33179;
			32358: outdata = 32'd33178;
			32359: outdata = 32'd33177;
			32360: outdata = 32'd33176;
			32361: outdata = 32'd33175;
			32362: outdata = 32'd33174;
			32363: outdata = 32'd33173;
			32364: outdata = 32'd33172;
			32365: outdata = 32'd33171;
			32366: outdata = 32'd33170;
			32367: outdata = 32'd33169;
			32368: outdata = 32'd33168;
			32369: outdata = 32'd33167;
			32370: outdata = 32'd33166;
			32371: outdata = 32'd33165;
			32372: outdata = 32'd33164;
			32373: outdata = 32'd33163;
			32374: outdata = 32'd33162;
			32375: outdata = 32'd33161;
			32376: outdata = 32'd33160;
			32377: outdata = 32'd33159;
			32378: outdata = 32'd33158;
			32379: outdata = 32'd33157;
			32380: outdata = 32'd33156;
			32381: outdata = 32'd33155;
			32382: outdata = 32'd33154;
			32383: outdata = 32'd33153;
			32384: outdata = 32'd33152;
			32385: outdata = 32'd33151;
			32386: outdata = 32'd33150;
			32387: outdata = 32'd33149;
			32388: outdata = 32'd33148;
			32389: outdata = 32'd33147;
			32390: outdata = 32'd33146;
			32391: outdata = 32'd33145;
			32392: outdata = 32'd33144;
			32393: outdata = 32'd33143;
			32394: outdata = 32'd33142;
			32395: outdata = 32'd33141;
			32396: outdata = 32'd33140;
			32397: outdata = 32'd33139;
			32398: outdata = 32'd33138;
			32399: outdata = 32'd33137;
			32400: outdata = 32'd33136;
			32401: outdata = 32'd33135;
			32402: outdata = 32'd33134;
			32403: outdata = 32'd33133;
			32404: outdata = 32'd33132;
			32405: outdata = 32'd33131;
			32406: outdata = 32'd33130;
			32407: outdata = 32'd33129;
			32408: outdata = 32'd33128;
			32409: outdata = 32'd33127;
			32410: outdata = 32'd33126;
			32411: outdata = 32'd33125;
			32412: outdata = 32'd33124;
			32413: outdata = 32'd33123;
			32414: outdata = 32'd33122;
			32415: outdata = 32'd33121;
			32416: outdata = 32'd33120;
			32417: outdata = 32'd33119;
			32418: outdata = 32'd33118;
			32419: outdata = 32'd33117;
			32420: outdata = 32'd33116;
			32421: outdata = 32'd33115;
			32422: outdata = 32'd33114;
			32423: outdata = 32'd33113;
			32424: outdata = 32'd33112;
			32425: outdata = 32'd33111;
			32426: outdata = 32'd33110;
			32427: outdata = 32'd33109;
			32428: outdata = 32'd33108;
			32429: outdata = 32'd33107;
			32430: outdata = 32'd33106;
			32431: outdata = 32'd33105;
			32432: outdata = 32'd33104;
			32433: outdata = 32'd33103;
			32434: outdata = 32'd33102;
			32435: outdata = 32'd33101;
			32436: outdata = 32'd33100;
			32437: outdata = 32'd33099;
			32438: outdata = 32'd33098;
			32439: outdata = 32'd33097;
			32440: outdata = 32'd33096;
			32441: outdata = 32'd33095;
			32442: outdata = 32'd33094;
			32443: outdata = 32'd33093;
			32444: outdata = 32'd33092;
			32445: outdata = 32'd33091;
			32446: outdata = 32'd33090;
			32447: outdata = 32'd33089;
			32448: outdata = 32'd33088;
			32449: outdata = 32'd33087;
			32450: outdata = 32'd33086;
			32451: outdata = 32'd33085;
			32452: outdata = 32'd33084;
			32453: outdata = 32'd33083;
			32454: outdata = 32'd33082;
			32455: outdata = 32'd33081;
			32456: outdata = 32'd33080;
			32457: outdata = 32'd33079;
			32458: outdata = 32'd33078;
			32459: outdata = 32'd33077;
			32460: outdata = 32'd33076;
			32461: outdata = 32'd33075;
			32462: outdata = 32'd33074;
			32463: outdata = 32'd33073;
			32464: outdata = 32'd33072;
			32465: outdata = 32'd33071;
			32466: outdata = 32'd33070;
			32467: outdata = 32'd33069;
			32468: outdata = 32'd33068;
			32469: outdata = 32'd33067;
			32470: outdata = 32'd33066;
			32471: outdata = 32'd33065;
			32472: outdata = 32'd33064;
			32473: outdata = 32'd33063;
			32474: outdata = 32'd33062;
			32475: outdata = 32'd33061;
			32476: outdata = 32'd33060;
			32477: outdata = 32'd33059;
			32478: outdata = 32'd33058;
			32479: outdata = 32'd33057;
			32480: outdata = 32'd33056;
			32481: outdata = 32'd33055;
			32482: outdata = 32'd33054;
			32483: outdata = 32'd33053;
			32484: outdata = 32'd33052;
			32485: outdata = 32'd33051;
			32486: outdata = 32'd33050;
			32487: outdata = 32'd33049;
			32488: outdata = 32'd33048;
			32489: outdata = 32'd33047;
			32490: outdata = 32'd33046;
			32491: outdata = 32'd33045;
			32492: outdata = 32'd33044;
			32493: outdata = 32'd33043;
			32494: outdata = 32'd33042;
			32495: outdata = 32'd33041;
			32496: outdata = 32'd33040;
			32497: outdata = 32'd33039;
			32498: outdata = 32'd33038;
			32499: outdata = 32'd33037;
			32500: outdata = 32'd33036;
			32501: outdata = 32'd33035;
			32502: outdata = 32'd33034;
			32503: outdata = 32'd33033;
			32504: outdata = 32'd33032;
			32505: outdata = 32'd33031;
			32506: outdata = 32'd33030;
			32507: outdata = 32'd33029;
			32508: outdata = 32'd33028;
			32509: outdata = 32'd33027;
			32510: outdata = 32'd33026;
			32511: outdata = 32'd33025;
			32512: outdata = 32'd33024;
			32513: outdata = 32'd33023;
			32514: outdata = 32'd33022;
			32515: outdata = 32'd33021;
			32516: outdata = 32'd33020;
			32517: outdata = 32'd33019;
			32518: outdata = 32'd33018;
			32519: outdata = 32'd33017;
			32520: outdata = 32'd33016;
			32521: outdata = 32'd33015;
			32522: outdata = 32'd33014;
			32523: outdata = 32'd33013;
			32524: outdata = 32'd33012;
			32525: outdata = 32'd33011;
			32526: outdata = 32'd33010;
			32527: outdata = 32'd33009;
			32528: outdata = 32'd33008;
			32529: outdata = 32'd33007;
			32530: outdata = 32'd33006;
			32531: outdata = 32'd33005;
			32532: outdata = 32'd33004;
			32533: outdata = 32'd33003;
			32534: outdata = 32'd33002;
			32535: outdata = 32'd33001;
			32536: outdata = 32'd33000;
			32537: outdata = 32'd32999;
			32538: outdata = 32'd32998;
			32539: outdata = 32'd32997;
			32540: outdata = 32'd32996;
			32541: outdata = 32'd32995;
			32542: outdata = 32'd32994;
			32543: outdata = 32'd32993;
			32544: outdata = 32'd32992;
			32545: outdata = 32'd32991;
			32546: outdata = 32'd32990;
			32547: outdata = 32'd32989;
			32548: outdata = 32'd32988;
			32549: outdata = 32'd32987;
			32550: outdata = 32'd32986;
			32551: outdata = 32'd32985;
			32552: outdata = 32'd32984;
			32553: outdata = 32'd32983;
			32554: outdata = 32'd32982;
			32555: outdata = 32'd32981;
			32556: outdata = 32'd32980;
			32557: outdata = 32'd32979;
			32558: outdata = 32'd32978;
			32559: outdata = 32'd32977;
			32560: outdata = 32'd32976;
			32561: outdata = 32'd32975;
			32562: outdata = 32'd32974;
			32563: outdata = 32'd32973;
			32564: outdata = 32'd32972;
			32565: outdata = 32'd32971;
			32566: outdata = 32'd32970;
			32567: outdata = 32'd32969;
			32568: outdata = 32'd32968;
			32569: outdata = 32'd32967;
			32570: outdata = 32'd32966;
			32571: outdata = 32'd32965;
			32572: outdata = 32'd32964;
			32573: outdata = 32'd32963;
			32574: outdata = 32'd32962;
			32575: outdata = 32'd32961;
			32576: outdata = 32'd32960;
			32577: outdata = 32'd32959;
			32578: outdata = 32'd32958;
			32579: outdata = 32'd32957;
			32580: outdata = 32'd32956;
			32581: outdata = 32'd32955;
			32582: outdata = 32'd32954;
			32583: outdata = 32'd32953;
			32584: outdata = 32'd32952;
			32585: outdata = 32'd32951;
			32586: outdata = 32'd32950;
			32587: outdata = 32'd32949;
			32588: outdata = 32'd32948;
			32589: outdata = 32'd32947;
			32590: outdata = 32'd32946;
			32591: outdata = 32'd32945;
			32592: outdata = 32'd32944;
			32593: outdata = 32'd32943;
			32594: outdata = 32'd32942;
			32595: outdata = 32'd32941;
			32596: outdata = 32'd32940;
			32597: outdata = 32'd32939;
			32598: outdata = 32'd32938;
			32599: outdata = 32'd32937;
			32600: outdata = 32'd32936;
			32601: outdata = 32'd32935;
			32602: outdata = 32'd32934;
			32603: outdata = 32'd32933;
			32604: outdata = 32'd32932;
			32605: outdata = 32'd32931;
			32606: outdata = 32'd32930;
			32607: outdata = 32'd32929;
			32608: outdata = 32'd32928;
			32609: outdata = 32'd32927;
			32610: outdata = 32'd32926;
			32611: outdata = 32'd32925;
			32612: outdata = 32'd32924;
			32613: outdata = 32'd32923;
			32614: outdata = 32'd32922;
			32615: outdata = 32'd32921;
			32616: outdata = 32'd32920;
			32617: outdata = 32'd32919;
			32618: outdata = 32'd32918;
			32619: outdata = 32'd32917;
			32620: outdata = 32'd32916;
			32621: outdata = 32'd32915;
			32622: outdata = 32'd32914;
			32623: outdata = 32'd32913;
			32624: outdata = 32'd32912;
			32625: outdata = 32'd32911;
			32626: outdata = 32'd32910;
			32627: outdata = 32'd32909;
			32628: outdata = 32'd32908;
			32629: outdata = 32'd32907;
			32630: outdata = 32'd32906;
			32631: outdata = 32'd32905;
			32632: outdata = 32'd32904;
			32633: outdata = 32'd32903;
			32634: outdata = 32'd32902;
			32635: outdata = 32'd32901;
			32636: outdata = 32'd32900;
			32637: outdata = 32'd32899;
			32638: outdata = 32'd32898;
			32639: outdata = 32'd32897;
			32640: outdata = 32'd32896;
			32641: outdata = 32'd32895;
			32642: outdata = 32'd32894;
			32643: outdata = 32'd32893;
			32644: outdata = 32'd32892;
			32645: outdata = 32'd32891;
			32646: outdata = 32'd32890;
			32647: outdata = 32'd32889;
			32648: outdata = 32'd32888;
			32649: outdata = 32'd32887;
			32650: outdata = 32'd32886;
			32651: outdata = 32'd32885;
			32652: outdata = 32'd32884;
			32653: outdata = 32'd32883;
			32654: outdata = 32'd32882;
			32655: outdata = 32'd32881;
			32656: outdata = 32'd32880;
			32657: outdata = 32'd32879;
			32658: outdata = 32'd32878;
			32659: outdata = 32'd32877;
			32660: outdata = 32'd32876;
			32661: outdata = 32'd32875;
			32662: outdata = 32'd32874;
			32663: outdata = 32'd32873;
			32664: outdata = 32'd32872;
			32665: outdata = 32'd32871;
			32666: outdata = 32'd32870;
			32667: outdata = 32'd32869;
			32668: outdata = 32'd32868;
			32669: outdata = 32'd32867;
			32670: outdata = 32'd32866;
			32671: outdata = 32'd32865;
			32672: outdata = 32'd32864;
			32673: outdata = 32'd32863;
			32674: outdata = 32'd32862;
			32675: outdata = 32'd32861;
			32676: outdata = 32'd32860;
			32677: outdata = 32'd32859;
			32678: outdata = 32'd32858;
			32679: outdata = 32'd32857;
			32680: outdata = 32'd32856;
			32681: outdata = 32'd32855;
			32682: outdata = 32'd32854;
			32683: outdata = 32'd32853;
			32684: outdata = 32'd32852;
			32685: outdata = 32'd32851;
			32686: outdata = 32'd32850;
			32687: outdata = 32'd32849;
			32688: outdata = 32'd32848;
			32689: outdata = 32'd32847;
			32690: outdata = 32'd32846;
			32691: outdata = 32'd32845;
			32692: outdata = 32'd32844;
			32693: outdata = 32'd32843;
			32694: outdata = 32'd32842;
			32695: outdata = 32'd32841;
			32696: outdata = 32'd32840;
			32697: outdata = 32'd32839;
			32698: outdata = 32'd32838;
			32699: outdata = 32'd32837;
			32700: outdata = 32'd32836;
			32701: outdata = 32'd32835;
			32702: outdata = 32'd32834;
			32703: outdata = 32'd32833;
			32704: outdata = 32'd32832;
			32705: outdata = 32'd32831;
			32706: outdata = 32'd32830;
			32707: outdata = 32'd32829;
			32708: outdata = 32'd32828;
			32709: outdata = 32'd32827;
			32710: outdata = 32'd32826;
			32711: outdata = 32'd32825;
			32712: outdata = 32'd32824;
			32713: outdata = 32'd32823;
			32714: outdata = 32'd32822;
			32715: outdata = 32'd32821;
			32716: outdata = 32'd32820;
			32717: outdata = 32'd32819;
			32718: outdata = 32'd32818;
			32719: outdata = 32'd32817;
			32720: outdata = 32'd32816;
			32721: outdata = 32'd32815;
			32722: outdata = 32'd32814;
			32723: outdata = 32'd32813;
			32724: outdata = 32'd32812;
			32725: outdata = 32'd32811;
			32726: outdata = 32'd32810;
			32727: outdata = 32'd32809;
			32728: outdata = 32'd32808;
			32729: outdata = 32'd32807;
			32730: outdata = 32'd32806;
			32731: outdata = 32'd32805;
			32732: outdata = 32'd32804;
			32733: outdata = 32'd32803;
			32734: outdata = 32'd32802;
			32735: outdata = 32'd32801;
			32736: outdata = 32'd32800;
			32737: outdata = 32'd32799;
			32738: outdata = 32'd32798;
			32739: outdata = 32'd32797;
			32740: outdata = 32'd32796;
			32741: outdata = 32'd32795;
			32742: outdata = 32'd32794;
			32743: outdata = 32'd32793;
			32744: outdata = 32'd32792;
			32745: outdata = 32'd32791;
			32746: outdata = 32'd32790;
			32747: outdata = 32'd32789;
			32748: outdata = 32'd32788;
			32749: outdata = 32'd32787;
			32750: outdata = 32'd32786;
			32751: outdata = 32'd32785;
			32752: outdata = 32'd32784;
			32753: outdata = 32'd32783;
			32754: outdata = 32'd32782;
			32755: outdata = 32'd32781;
			32756: outdata = 32'd32780;
			32757: outdata = 32'd32779;
			32758: outdata = 32'd32778;
			32759: outdata = 32'd32777;
			32760: outdata = 32'd32776;
			32761: outdata = 32'd32775;
			32762: outdata = 32'd32774;
			32763: outdata = 32'd32773;
			32764: outdata = 32'd32772;
			32765: outdata = 32'd32771;
			32766: outdata = 32'd32770;
			32767: outdata = 32'd32769;
			32768: outdata = 32'd32768;
			32769: outdata = 32'd32767;
			32770: outdata = 32'd32766;
			32771: outdata = 32'd32765;
			32772: outdata = 32'd32764;
			32773: outdata = 32'd32763;
			32774: outdata = 32'd32762;
			32775: outdata = 32'd32761;
			32776: outdata = 32'd32760;
			32777: outdata = 32'd32759;
			32778: outdata = 32'd32758;
			32779: outdata = 32'd32757;
			32780: outdata = 32'd32756;
			32781: outdata = 32'd32755;
			32782: outdata = 32'd32754;
			32783: outdata = 32'd32753;
			32784: outdata = 32'd32752;
			32785: outdata = 32'd32751;
			32786: outdata = 32'd32750;
			32787: outdata = 32'd32749;
			32788: outdata = 32'd32748;
			32789: outdata = 32'd32747;
			32790: outdata = 32'd32746;
			32791: outdata = 32'd32745;
			32792: outdata = 32'd32744;
			32793: outdata = 32'd32743;
			32794: outdata = 32'd32742;
			32795: outdata = 32'd32741;
			32796: outdata = 32'd32740;
			32797: outdata = 32'd32739;
			32798: outdata = 32'd32738;
			32799: outdata = 32'd32737;
			32800: outdata = 32'd32736;
			32801: outdata = 32'd32735;
			32802: outdata = 32'd32734;
			32803: outdata = 32'd32733;
			32804: outdata = 32'd32732;
			32805: outdata = 32'd32731;
			32806: outdata = 32'd32730;
			32807: outdata = 32'd32729;
			32808: outdata = 32'd32728;
			32809: outdata = 32'd32727;
			32810: outdata = 32'd32726;
			32811: outdata = 32'd32725;
			32812: outdata = 32'd32724;
			32813: outdata = 32'd32723;
			32814: outdata = 32'd32722;
			32815: outdata = 32'd32721;
			32816: outdata = 32'd32720;
			32817: outdata = 32'd32719;
			32818: outdata = 32'd32718;
			32819: outdata = 32'd32717;
			32820: outdata = 32'd32716;
			32821: outdata = 32'd32715;
			32822: outdata = 32'd32714;
			32823: outdata = 32'd32713;
			32824: outdata = 32'd32712;
			32825: outdata = 32'd32711;
			32826: outdata = 32'd32710;
			32827: outdata = 32'd32709;
			32828: outdata = 32'd32708;
			32829: outdata = 32'd32707;
			32830: outdata = 32'd32706;
			32831: outdata = 32'd32705;
			32832: outdata = 32'd32704;
			32833: outdata = 32'd32703;
			32834: outdata = 32'd32702;
			32835: outdata = 32'd32701;
			32836: outdata = 32'd32700;
			32837: outdata = 32'd32699;
			32838: outdata = 32'd32698;
			32839: outdata = 32'd32697;
			32840: outdata = 32'd32696;
			32841: outdata = 32'd32695;
			32842: outdata = 32'd32694;
			32843: outdata = 32'd32693;
			32844: outdata = 32'd32692;
			32845: outdata = 32'd32691;
			32846: outdata = 32'd32690;
			32847: outdata = 32'd32689;
			32848: outdata = 32'd32688;
			32849: outdata = 32'd32687;
			32850: outdata = 32'd32686;
			32851: outdata = 32'd32685;
			32852: outdata = 32'd32684;
			32853: outdata = 32'd32683;
			32854: outdata = 32'd32682;
			32855: outdata = 32'd32681;
			32856: outdata = 32'd32680;
			32857: outdata = 32'd32679;
			32858: outdata = 32'd32678;
			32859: outdata = 32'd32677;
			32860: outdata = 32'd32676;
			32861: outdata = 32'd32675;
			32862: outdata = 32'd32674;
			32863: outdata = 32'd32673;
			32864: outdata = 32'd32672;
			32865: outdata = 32'd32671;
			32866: outdata = 32'd32670;
			32867: outdata = 32'd32669;
			32868: outdata = 32'd32668;
			32869: outdata = 32'd32667;
			32870: outdata = 32'd32666;
			32871: outdata = 32'd32665;
			32872: outdata = 32'd32664;
			32873: outdata = 32'd32663;
			32874: outdata = 32'd32662;
			32875: outdata = 32'd32661;
			32876: outdata = 32'd32660;
			32877: outdata = 32'd32659;
			32878: outdata = 32'd32658;
			32879: outdata = 32'd32657;
			32880: outdata = 32'd32656;
			32881: outdata = 32'd32655;
			32882: outdata = 32'd32654;
			32883: outdata = 32'd32653;
			32884: outdata = 32'd32652;
			32885: outdata = 32'd32651;
			32886: outdata = 32'd32650;
			32887: outdata = 32'd32649;
			32888: outdata = 32'd32648;
			32889: outdata = 32'd32647;
			32890: outdata = 32'd32646;
			32891: outdata = 32'd32645;
			32892: outdata = 32'd32644;
			32893: outdata = 32'd32643;
			32894: outdata = 32'd32642;
			32895: outdata = 32'd32641;
			32896: outdata = 32'd32640;
			32897: outdata = 32'd32639;
			32898: outdata = 32'd32638;
			32899: outdata = 32'd32637;
			32900: outdata = 32'd32636;
			32901: outdata = 32'd32635;
			32902: outdata = 32'd32634;
			32903: outdata = 32'd32633;
			32904: outdata = 32'd32632;
			32905: outdata = 32'd32631;
			32906: outdata = 32'd32630;
			32907: outdata = 32'd32629;
			32908: outdata = 32'd32628;
			32909: outdata = 32'd32627;
			32910: outdata = 32'd32626;
			32911: outdata = 32'd32625;
			32912: outdata = 32'd32624;
			32913: outdata = 32'd32623;
			32914: outdata = 32'd32622;
			32915: outdata = 32'd32621;
			32916: outdata = 32'd32620;
			32917: outdata = 32'd32619;
			32918: outdata = 32'd32618;
			32919: outdata = 32'd32617;
			32920: outdata = 32'd32616;
			32921: outdata = 32'd32615;
			32922: outdata = 32'd32614;
			32923: outdata = 32'd32613;
			32924: outdata = 32'd32612;
			32925: outdata = 32'd32611;
			32926: outdata = 32'd32610;
			32927: outdata = 32'd32609;
			32928: outdata = 32'd32608;
			32929: outdata = 32'd32607;
			32930: outdata = 32'd32606;
			32931: outdata = 32'd32605;
			32932: outdata = 32'd32604;
			32933: outdata = 32'd32603;
			32934: outdata = 32'd32602;
			32935: outdata = 32'd32601;
			32936: outdata = 32'd32600;
			32937: outdata = 32'd32599;
			32938: outdata = 32'd32598;
			32939: outdata = 32'd32597;
			32940: outdata = 32'd32596;
			32941: outdata = 32'd32595;
			32942: outdata = 32'd32594;
			32943: outdata = 32'd32593;
			32944: outdata = 32'd32592;
			32945: outdata = 32'd32591;
			32946: outdata = 32'd32590;
			32947: outdata = 32'd32589;
			32948: outdata = 32'd32588;
			32949: outdata = 32'd32587;
			32950: outdata = 32'd32586;
			32951: outdata = 32'd32585;
			32952: outdata = 32'd32584;
			32953: outdata = 32'd32583;
			32954: outdata = 32'd32582;
			32955: outdata = 32'd32581;
			32956: outdata = 32'd32580;
			32957: outdata = 32'd32579;
			32958: outdata = 32'd32578;
			32959: outdata = 32'd32577;
			32960: outdata = 32'd32576;
			32961: outdata = 32'd32575;
			32962: outdata = 32'd32574;
			32963: outdata = 32'd32573;
			32964: outdata = 32'd32572;
			32965: outdata = 32'd32571;
			32966: outdata = 32'd32570;
			32967: outdata = 32'd32569;
			32968: outdata = 32'd32568;
			32969: outdata = 32'd32567;
			32970: outdata = 32'd32566;
			32971: outdata = 32'd32565;
			32972: outdata = 32'd32564;
			32973: outdata = 32'd32563;
			32974: outdata = 32'd32562;
			32975: outdata = 32'd32561;
			32976: outdata = 32'd32560;
			32977: outdata = 32'd32559;
			32978: outdata = 32'd32558;
			32979: outdata = 32'd32557;
			32980: outdata = 32'd32556;
			32981: outdata = 32'd32555;
			32982: outdata = 32'd32554;
			32983: outdata = 32'd32553;
			32984: outdata = 32'd32552;
			32985: outdata = 32'd32551;
			32986: outdata = 32'd32550;
			32987: outdata = 32'd32549;
			32988: outdata = 32'd32548;
			32989: outdata = 32'd32547;
			32990: outdata = 32'd32546;
			32991: outdata = 32'd32545;
			32992: outdata = 32'd32544;
			32993: outdata = 32'd32543;
			32994: outdata = 32'd32542;
			32995: outdata = 32'd32541;
			32996: outdata = 32'd32540;
			32997: outdata = 32'd32539;
			32998: outdata = 32'd32538;
			32999: outdata = 32'd32537;
			33000: outdata = 32'd32536;
			33001: outdata = 32'd32535;
			33002: outdata = 32'd32534;
			33003: outdata = 32'd32533;
			33004: outdata = 32'd32532;
			33005: outdata = 32'd32531;
			33006: outdata = 32'd32530;
			33007: outdata = 32'd32529;
			33008: outdata = 32'd32528;
			33009: outdata = 32'd32527;
			33010: outdata = 32'd32526;
			33011: outdata = 32'd32525;
			33012: outdata = 32'd32524;
			33013: outdata = 32'd32523;
			33014: outdata = 32'd32522;
			33015: outdata = 32'd32521;
			33016: outdata = 32'd32520;
			33017: outdata = 32'd32519;
			33018: outdata = 32'd32518;
			33019: outdata = 32'd32517;
			33020: outdata = 32'd32516;
			33021: outdata = 32'd32515;
			33022: outdata = 32'd32514;
			33023: outdata = 32'd32513;
			33024: outdata = 32'd32512;
			33025: outdata = 32'd32511;
			33026: outdata = 32'd32510;
			33027: outdata = 32'd32509;
			33028: outdata = 32'd32508;
			33029: outdata = 32'd32507;
			33030: outdata = 32'd32506;
			33031: outdata = 32'd32505;
			33032: outdata = 32'd32504;
			33033: outdata = 32'd32503;
			33034: outdata = 32'd32502;
			33035: outdata = 32'd32501;
			33036: outdata = 32'd32500;
			33037: outdata = 32'd32499;
			33038: outdata = 32'd32498;
			33039: outdata = 32'd32497;
			33040: outdata = 32'd32496;
			33041: outdata = 32'd32495;
			33042: outdata = 32'd32494;
			33043: outdata = 32'd32493;
			33044: outdata = 32'd32492;
			33045: outdata = 32'd32491;
			33046: outdata = 32'd32490;
			33047: outdata = 32'd32489;
			33048: outdata = 32'd32488;
			33049: outdata = 32'd32487;
			33050: outdata = 32'd32486;
			33051: outdata = 32'd32485;
			33052: outdata = 32'd32484;
			33053: outdata = 32'd32483;
			33054: outdata = 32'd32482;
			33055: outdata = 32'd32481;
			33056: outdata = 32'd32480;
			33057: outdata = 32'd32479;
			33058: outdata = 32'd32478;
			33059: outdata = 32'd32477;
			33060: outdata = 32'd32476;
			33061: outdata = 32'd32475;
			33062: outdata = 32'd32474;
			33063: outdata = 32'd32473;
			33064: outdata = 32'd32472;
			33065: outdata = 32'd32471;
			33066: outdata = 32'd32470;
			33067: outdata = 32'd32469;
			33068: outdata = 32'd32468;
			33069: outdata = 32'd32467;
			33070: outdata = 32'd32466;
			33071: outdata = 32'd32465;
			33072: outdata = 32'd32464;
			33073: outdata = 32'd32463;
			33074: outdata = 32'd32462;
			33075: outdata = 32'd32461;
			33076: outdata = 32'd32460;
			33077: outdata = 32'd32459;
			33078: outdata = 32'd32458;
			33079: outdata = 32'd32457;
			33080: outdata = 32'd32456;
			33081: outdata = 32'd32455;
			33082: outdata = 32'd32454;
			33083: outdata = 32'd32453;
			33084: outdata = 32'd32452;
			33085: outdata = 32'd32451;
			33086: outdata = 32'd32450;
			33087: outdata = 32'd32449;
			33088: outdata = 32'd32448;
			33089: outdata = 32'd32447;
			33090: outdata = 32'd32446;
			33091: outdata = 32'd32445;
			33092: outdata = 32'd32444;
			33093: outdata = 32'd32443;
			33094: outdata = 32'd32442;
			33095: outdata = 32'd32441;
			33096: outdata = 32'd32440;
			33097: outdata = 32'd32439;
			33098: outdata = 32'd32438;
			33099: outdata = 32'd32437;
			33100: outdata = 32'd32436;
			33101: outdata = 32'd32435;
			33102: outdata = 32'd32434;
			33103: outdata = 32'd32433;
			33104: outdata = 32'd32432;
			33105: outdata = 32'd32431;
			33106: outdata = 32'd32430;
			33107: outdata = 32'd32429;
			33108: outdata = 32'd32428;
			33109: outdata = 32'd32427;
			33110: outdata = 32'd32426;
			33111: outdata = 32'd32425;
			33112: outdata = 32'd32424;
			33113: outdata = 32'd32423;
			33114: outdata = 32'd32422;
			33115: outdata = 32'd32421;
			33116: outdata = 32'd32420;
			33117: outdata = 32'd32419;
			33118: outdata = 32'd32418;
			33119: outdata = 32'd32417;
			33120: outdata = 32'd32416;
			33121: outdata = 32'd32415;
			33122: outdata = 32'd32414;
			33123: outdata = 32'd32413;
			33124: outdata = 32'd32412;
			33125: outdata = 32'd32411;
			33126: outdata = 32'd32410;
			33127: outdata = 32'd32409;
			33128: outdata = 32'd32408;
			33129: outdata = 32'd32407;
			33130: outdata = 32'd32406;
			33131: outdata = 32'd32405;
			33132: outdata = 32'd32404;
			33133: outdata = 32'd32403;
			33134: outdata = 32'd32402;
			33135: outdata = 32'd32401;
			33136: outdata = 32'd32400;
			33137: outdata = 32'd32399;
			33138: outdata = 32'd32398;
			33139: outdata = 32'd32397;
			33140: outdata = 32'd32396;
			33141: outdata = 32'd32395;
			33142: outdata = 32'd32394;
			33143: outdata = 32'd32393;
			33144: outdata = 32'd32392;
			33145: outdata = 32'd32391;
			33146: outdata = 32'd32390;
			33147: outdata = 32'd32389;
			33148: outdata = 32'd32388;
			33149: outdata = 32'd32387;
			33150: outdata = 32'd32386;
			33151: outdata = 32'd32385;
			33152: outdata = 32'd32384;
			33153: outdata = 32'd32383;
			33154: outdata = 32'd32382;
			33155: outdata = 32'd32381;
			33156: outdata = 32'd32380;
			33157: outdata = 32'd32379;
			33158: outdata = 32'd32378;
			33159: outdata = 32'd32377;
			33160: outdata = 32'd32376;
			33161: outdata = 32'd32375;
			33162: outdata = 32'd32374;
			33163: outdata = 32'd32373;
			33164: outdata = 32'd32372;
			33165: outdata = 32'd32371;
			33166: outdata = 32'd32370;
			33167: outdata = 32'd32369;
			33168: outdata = 32'd32368;
			33169: outdata = 32'd32367;
			33170: outdata = 32'd32366;
			33171: outdata = 32'd32365;
			33172: outdata = 32'd32364;
			33173: outdata = 32'd32363;
			33174: outdata = 32'd32362;
			33175: outdata = 32'd32361;
			33176: outdata = 32'd32360;
			33177: outdata = 32'd32359;
			33178: outdata = 32'd32358;
			33179: outdata = 32'd32357;
			33180: outdata = 32'd32356;
			33181: outdata = 32'd32355;
			33182: outdata = 32'd32354;
			33183: outdata = 32'd32353;
			33184: outdata = 32'd32352;
			33185: outdata = 32'd32351;
			33186: outdata = 32'd32350;
			33187: outdata = 32'd32349;
			33188: outdata = 32'd32348;
			33189: outdata = 32'd32347;
			33190: outdata = 32'd32346;
			33191: outdata = 32'd32345;
			33192: outdata = 32'd32344;
			33193: outdata = 32'd32343;
			33194: outdata = 32'd32342;
			33195: outdata = 32'd32341;
			33196: outdata = 32'd32340;
			33197: outdata = 32'd32339;
			33198: outdata = 32'd32338;
			33199: outdata = 32'd32337;
			33200: outdata = 32'd32336;
			33201: outdata = 32'd32335;
			33202: outdata = 32'd32334;
			33203: outdata = 32'd32333;
			33204: outdata = 32'd32332;
			33205: outdata = 32'd32331;
			33206: outdata = 32'd32330;
			33207: outdata = 32'd32329;
			33208: outdata = 32'd32328;
			33209: outdata = 32'd32327;
			33210: outdata = 32'd32326;
			33211: outdata = 32'd32325;
			33212: outdata = 32'd32324;
			33213: outdata = 32'd32323;
			33214: outdata = 32'd32322;
			33215: outdata = 32'd32321;
			33216: outdata = 32'd32320;
			33217: outdata = 32'd32319;
			33218: outdata = 32'd32318;
			33219: outdata = 32'd32317;
			33220: outdata = 32'd32316;
			33221: outdata = 32'd32315;
			33222: outdata = 32'd32314;
			33223: outdata = 32'd32313;
			33224: outdata = 32'd32312;
			33225: outdata = 32'd32311;
			33226: outdata = 32'd32310;
			33227: outdata = 32'd32309;
			33228: outdata = 32'd32308;
			33229: outdata = 32'd32307;
			33230: outdata = 32'd32306;
			33231: outdata = 32'd32305;
			33232: outdata = 32'd32304;
			33233: outdata = 32'd32303;
			33234: outdata = 32'd32302;
			33235: outdata = 32'd32301;
			33236: outdata = 32'd32300;
			33237: outdata = 32'd32299;
			33238: outdata = 32'd32298;
			33239: outdata = 32'd32297;
			33240: outdata = 32'd32296;
			33241: outdata = 32'd32295;
			33242: outdata = 32'd32294;
			33243: outdata = 32'd32293;
			33244: outdata = 32'd32292;
			33245: outdata = 32'd32291;
			33246: outdata = 32'd32290;
			33247: outdata = 32'd32289;
			33248: outdata = 32'd32288;
			33249: outdata = 32'd32287;
			33250: outdata = 32'd32286;
			33251: outdata = 32'd32285;
			33252: outdata = 32'd32284;
			33253: outdata = 32'd32283;
			33254: outdata = 32'd32282;
			33255: outdata = 32'd32281;
			33256: outdata = 32'd32280;
			33257: outdata = 32'd32279;
			33258: outdata = 32'd32278;
			33259: outdata = 32'd32277;
			33260: outdata = 32'd32276;
			33261: outdata = 32'd32275;
			33262: outdata = 32'd32274;
			33263: outdata = 32'd32273;
			33264: outdata = 32'd32272;
			33265: outdata = 32'd32271;
			33266: outdata = 32'd32270;
			33267: outdata = 32'd32269;
			33268: outdata = 32'd32268;
			33269: outdata = 32'd32267;
			33270: outdata = 32'd32266;
			33271: outdata = 32'd32265;
			33272: outdata = 32'd32264;
			33273: outdata = 32'd32263;
			33274: outdata = 32'd32262;
			33275: outdata = 32'd32261;
			33276: outdata = 32'd32260;
			33277: outdata = 32'd32259;
			33278: outdata = 32'd32258;
			33279: outdata = 32'd32257;
			33280: outdata = 32'd32256;
			33281: outdata = 32'd32255;
			33282: outdata = 32'd32254;
			33283: outdata = 32'd32253;
			33284: outdata = 32'd32252;
			33285: outdata = 32'd32251;
			33286: outdata = 32'd32250;
			33287: outdata = 32'd32249;
			33288: outdata = 32'd32248;
			33289: outdata = 32'd32247;
			33290: outdata = 32'd32246;
			33291: outdata = 32'd32245;
			33292: outdata = 32'd32244;
			33293: outdata = 32'd32243;
			33294: outdata = 32'd32242;
			33295: outdata = 32'd32241;
			33296: outdata = 32'd32240;
			33297: outdata = 32'd32239;
			33298: outdata = 32'd32238;
			33299: outdata = 32'd32237;
			33300: outdata = 32'd32236;
			33301: outdata = 32'd32235;
			33302: outdata = 32'd32234;
			33303: outdata = 32'd32233;
			33304: outdata = 32'd32232;
			33305: outdata = 32'd32231;
			33306: outdata = 32'd32230;
			33307: outdata = 32'd32229;
			33308: outdata = 32'd32228;
			33309: outdata = 32'd32227;
			33310: outdata = 32'd32226;
			33311: outdata = 32'd32225;
			33312: outdata = 32'd32224;
			33313: outdata = 32'd32223;
			33314: outdata = 32'd32222;
			33315: outdata = 32'd32221;
			33316: outdata = 32'd32220;
			33317: outdata = 32'd32219;
			33318: outdata = 32'd32218;
			33319: outdata = 32'd32217;
			33320: outdata = 32'd32216;
			33321: outdata = 32'd32215;
			33322: outdata = 32'd32214;
			33323: outdata = 32'd32213;
			33324: outdata = 32'd32212;
			33325: outdata = 32'd32211;
			33326: outdata = 32'd32210;
			33327: outdata = 32'd32209;
			33328: outdata = 32'd32208;
			33329: outdata = 32'd32207;
			33330: outdata = 32'd32206;
			33331: outdata = 32'd32205;
			33332: outdata = 32'd32204;
			33333: outdata = 32'd32203;
			33334: outdata = 32'd32202;
			33335: outdata = 32'd32201;
			33336: outdata = 32'd32200;
			33337: outdata = 32'd32199;
			33338: outdata = 32'd32198;
			33339: outdata = 32'd32197;
			33340: outdata = 32'd32196;
			33341: outdata = 32'd32195;
			33342: outdata = 32'd32194;
			33343: outdata = 32'd32193;
			33344: outdata = 32'd32192;
			33345: outdata = 32'd32191;
			33346: outdata = 32'd32190;
			33347: outdata = 32'd32189;
			33348: outdata = 32'd32188;
			33349: outdata = 32'd32187;
			33350: outdata = 32'd32186;
			33351: outdata = 32'd32185;
			33352: outdata = 32'd32184;
			33353: outdata = 32'd32183;
			33354: outdata = 32'd32182;
			33355: outdata = 32'd32181;
			33356: outdata = 32'd32180;
			33357: outdata = 32'd32179;
			33358: outdata = 32'd32178;
			33359: outdata = 32'd32177;
			33360: outdata = 32'd32176;
			33361: outdata = 32'd32175;
			33362: outdata = 32'd32174;
			33363: outdata = 32'd32173;
			33364: outdata = 32'd32172;
			33365: outdata = 32'd32171;
			33366: outdata = 32'd32170;
			33367: outdata = 32'd32169;
			33368: outdata = 32'd32168;
			33369: outdata = 32'd32167;
			33370: outdata = 32'd32166;
			33371: outdata = 32'd32165;
			33372: outdata = 32'd32164;
			33373: outdata = 32'd32163;
			33374: outdata = 32'd32162;
			33375: outdata = 32'd32161;
			33376: outdata = 32'd32160;
			33377: outdata = 32'd32159;
			33378: outdata = 32'd32158;
			33379: outdata = 32'd32157;
			33380: outdata = 32'd32156;
			33381: outdata = 32'd32155;
			33382: outdata = 32'd32154;
			33383: outdata = 32'd32153;
			33384: outdata = 32'd32152;
			33385: outdata = 32'd32151;
			33386: outdata = 32'd32150;
			33387: outdata = 32'd32149;
			33388: outdata = 32'd32148;
			33389: outdata = 32'd32147;
			33390: outdata = 32'd32146;
			33391: outdata = 32'd32145;
			33392: outdata = 32'd32144;
			33393: outdata = 32'd32143;
			33394: outdata = 32'd32142;
			33395: outdata = 32'd32141;
			33396: outdata = 32'd32140;
			33397: outdata = 32'd32139;
			33398: outdata = 32'd32138;
			33399: outdata = 32'd32137;
			33400: outdata = 32'd32136;
			33401: outdata = 32'd32135;
			33402: outdata = 32'd32134;
			33403: outdata = 32'd32133;
			33404: outdata = 32'd32132;
			33405: outdata = 32'd32131;
			33406: outdata = 32'd32130;
			33407: outdata = 32'd32129;
			33408: outdata = 32'd32128;
			33409: outdata = 32'd32127;
			33410: outdata = 32'd32126;
			33411: outdata = 32'd32125;
			33412: outdata = 32'd32124;
			33413: outdata = 32'd32123;
			33414: outdata = 32'd32122;
			33415: outdata = 32'd32121;
			33416: outdata = 32'd32120;
			33417: outdata = 32'd32119;
			33418: outdata = 32'd32118;
			33419: outdata = 32'd32117;
			33420: outdata = 32'd32116;
			33421: outdata = 32'd32115;
			33422: outdata = 32'd32114;
			33423: outdata = 32'd32113;
			33424: outdata = 32'd32112;
			33425: outdata = 32'd32111;
			33426: outdata = 32'd32110;
			33427: outdata = 32'd32109;
			33428: outdata = 32'd32108;
			33429: outdata = 32'd32107;
			33430: outdata = 32'd32106;
			33431: outdata = 32'd32105;
			33432: outdata = 32'd32104;
			33433: outdata = 32'd32103;
			33434: outdata = 32'd32102;
			33435: outdata = 32'd32101;
			33436: outdata = 32'd32100;
			33437: outdata = 32'd32099;
			33438: outdata = 32'd32098;
			33439: outdata = 32'd32097;
			33440: outdata = 32'd32096;
			33441: outdata = 32'd32095;
			33442: outdata = 32'd32094;
			33443: outdata = 32'd32093;
			33444: outdata = 32'd32092;
			33445: outdata = 32'd32091;
			33446: outdata = 32'd32090;
			33447: outdata = 32'd32089;
			33448: outdata = 32'd32088;
			33449: outdata = 32'd32087;
			33450: outdata = 32'd32086;
			33451: outdata = 32'd32085;
			33452: outdata = 32'd32084;
			33453: outdata = 32'd32083;
			33454: outdata = 32'd32082;
			33455: outdata = 32'd32081;
			33456: outdata = 32'd32080;
			33457: outdata = 32'd32079;
			33458: outdata = 32'd32078;
			33459: outdata = 32'd32077;
			33460: outdata = 32'd32076;
			33461: outdata = 32'd32075;
			33462: outdata = 32'd32074;
			33463: outdata = 32'd32073;
			33464: outdata = 32'd32072;
			33465: outdata = 32'd32071;
			33466: outdata = 32'd32070;
			33467: outdata = 32'd32069;
			33468: outdata = 32'd32068;
			33469: outdata = 32'd32067;
			33470: outdata = 32'd32066;
			33471: outdata = 32'd32065;
			33472: outdata = 32'd32064;
			33473: outdata = 32'd32063;
			33474: outdata = 32'd32062;
			33475: outdata = 32'd32061;
			33476: outdata = 32'd32060;
			33477: outdata = 32'd32059;
			33478: outdata = 32'd32058;
			33479: outdata = 32'd32057;
			33480: outdata = 32'd32056;
			33481: outdata = 32'd32055;
			33482: outdata = 32'd32054;
			33483: outdata = 32'd32053;
			33484: outdata = 32'd32052;
			33485: outdata = 32'd32051;
			33486: outdata = 32'd32050;
			33487: outdata = 32'd32049;
			33488: outdata = 32'd32048;
			33489: outdata = 32'd32047;
			33490: outdata = 32'd32046;
			33491: outdata = 32'd32045;
			33492: outdata = 32'd32044;
			33493: outdata = 32'd32043;
			33494: outdata = 32'd32042;
			33495: outdata = 32'd32041;
			33496: outdata = 32'd32040;
			33497: outdata = 32'd32039;
			33498: outdata = 32'd32038;
			33499: outdata = 32'd32037;
			33500: outdata = 32'd32036;
			33501: outdata = 32'd32035;
			33502: outdata = 32'd32034;
			33503: outdata = 32'd32033;
			33504: outdata = 32'd32032;
			33505: outdata = 32'd32031;
			33506: outdata = 32'd32030;
			33507: outdata = 32'd32029;
			33508: outdata = 32'd32028;
			33509: outdata = 32'd32027;
			33510: outdata = 32'd32026;
			33511: outdata = 32'd32025;
			33512: outdata = 32'd32024;
			33513: outdata = 32'd32023;
			33514: outdata = 32'd32022;
			33515: outdata = 32'd32021;
			33516: outdata = 32'd32020;
			33517: outdata = 32'd32019;
			33518: outdata = 32'd32018;
			33519: outdata = 32'd32017;
			33520: outdata = 32'd32016;
			33521: outdata = 32'd32015;
			33522: outdata = 32'd32014;
			33523: outdata = 32'd32013;
			33524: outdata = 32'd32012;
			33525: outdata = 32'd32011;
			33526: outdata = 32'd32010;
			33527: outdata = 32'd32009;
			33528: outdata = 32'd32008;
			33529: outdata = 32'd32007;
			33530: outdata = 32'd32006;
			33531: outdata = 32'd32005;
			33532: outdata = 32'd32004;
			33533: outdata = 32'd32003;
			33534: outdata = 32'd32002;
			33535: outdata = 32'd32001;
			33536: outdata = 32'd32000;
			33537: outdata = 32'd31999;
			33538: outdata = 32'd31998;
			33539: outdata = 32'd31997;
			33540: outdata = 32'd31996;
			33541: outdata = 32'd31995;
			33542: outdata = 32'd31994;
			33543: outdata = 32'd31993;
			33544: outdata = 32'd31992;
			33545: outdata = 32'd31991;
			33546: outdata = 32'd31990;
			33547: outdata = 32'd31989;
			33548: outdata = 32'd31988;
			33549: outdata = 32'd31987;
			33550: outdata = 32'd31986;
			33551: outdata = 32'd31985;
			33552: outdata = 32'd31984;
			33553: outdata = 32'd31983;
			33554: outdata = 32'd31982;
			33555: outdata = 32'd31981;
			33556: outdata = 32'd31980;
			33557: outdata = 32'd31979;
			33558: outdata = 32'd31978;
			33559: outdata = 32'd31977;
			33560: outdata = 32'd31976;
			33561: outdata = 32'd31975;
			33562: outdata = 32'd31974;
			33563: outdata = 32'd31973;
			33564: outdata = 32'd31972;
			33565: outdata = 32'd31971;
			33566: outdata = 32'd31970;
			33567: outdata = 32'd31969;
			33568: outdata = 32'd31968;
			33569: outdata = 32'd31967;
			33570: outdata = 32'd31966;
			33571: outdata = 32'd31965;
			33572: outdata = 32'd31964;
			33573: outdata = 32'd31963;
			33574: outdata = 32'd31962;
			33575: outdata = 32'd31961;
			33576: outdata = 32'd31960;
			33577: outdata = 32'd31959;
			33578: outdata = 32'd31958;
			33579: outdata = 32'd31957;
			33580: outdata = 32'd31956;
			33581: outdata = 32'd31955;
			33582: outdata = 32'd31954;
			33583: outdata = 32'd31953;
			33584: outdata = 32'd31952;
			33585: outdata = 32'd31951;
			33586: outdata = 32'd31950;
			33587: outdata = 32'd31949;
			33588: outdata = 32'd31948;
			33589: outdata = 32'd31947;
			33590: outdata = 32'd31946;
			33591: outdata = 32'd31945;
			33592: outdata = 32'd31944;
			33593: outdata = 32'd31943;
			33594: outdata = 32'd31942;
			33595: outdata = 32'd31941;
			33596: outdata = 32'd31940;
			33597: outdata = 32'd31939;
			33598: outdata = 32'd31938;
			33599: outdata = 32'd31937;
			33600: outdata = 32'd31936;
			33601: outdata = 32'd31935;
			33602: outdata = 32'd31934;
			33603: outdata = 32'd31933;
			33604: outdata = 32'd31932;
			33605: outdata = 32'd31931;
			33606: outdata = 32'd31930;
			33607: outdata = 32'd31929;
			33608: outdata = 32'd31928;
			33609: outdata = 32'd31927;
			33610: outdata = 32'd31926;
			33611: outdata = 32'd31925;
			33612: outdata = 32'd31924;
			33613: outdata = 32'd31923;
			33614: outdata = 32'd31922;
			33615: outdata = 32'd31921;
			33616: outdata = 32'd31920;
			33617: outdata = 32'd31919;
			33618: outdata = 32'd31918;
			33619: outdata = 32'd31917;
			33620: outdata = 32'd31916;
			33621: outdata = 32'd31915;
			33622: outdata = 32'd31914;
			33623: outdata = 32'd31913;
			33624: outdata = 32'd31912;
			33625: outdata = 32'd31911;
			33626: outdata = 32'd31910;
			33627: outdata = 32'd31909;
			33628: outdata = 32'd31908;
			33629: outdata = 32'd31907;
			33630: outdata = 32'd31906;
			33631: outdata = 32'd31905;
			33632: outdata = 32'd31904;
			33633: outdata = 32'd31903;
			33634: outdata = 32'd31902;
			33635: outdata = 32'd31901;
			33636: outdata = 32'd31900;
			33637: outdata = 32'd31899;
			33638: outdata = 32'd31898;
			33639: outdata = 32'd31897;
			33640: outdata = 32'd31896;
			33641: outdata = 32'd31895;
			33642: outdata = 32'd31894;
			33643: outdata = 32'd31893;
			33644: outdata = 32'd31892;
			33645: outdata = 32'd31891;
			33646: outdata = 32'd31890;
			33647: outdata = 32'd31889;
			33648: outdata = 32'd31888;
			33649: outdata = 32'd31887;
			33650: outdata = 32'd31886;
			33651: outdata = 32'd31885;
			33652: outdata = 32'd31884;
			33653: outdata = 32'd31883;
			33654: outdata = 32'd31882;
			33655: outdata = 32'd31881;
			33656: outdata = 32'd31880;
			33657: outdata = 32'd31879;
			33658: outdata = 32'd31878;
			33659: outdata = 32'd31877;
			33660: outdata = 32'd31876;
			33661: outdata = 32'd31875;
			33662: outdata = 32'd31874;
			33663: outdata = 32'd31873;
			33664: outdata = 32'd31872;
			33665: outdata = 32'd31871;
			33666: outdata = 32'd31870;
			33667: outdata = 32'd31869;
			33668: outdata = 32'd31868;
			33669: outdata = 32'd31867;
			33670: outdata = 32'd31866;
			33671: outdata = 32'd31865;
			33672: outdata = 32'd31864;
			33673: outdata = 32'd31863;
			33674: outdata = 32'd31862;
			33675: outdata = 32'd31861;
			33676: outdata = 32'd31860;
			33677: outdata = 32'd31859;
			33678: outdata = 32'd31858;
			33679: outdata = 32'd31857;
			33680: outdata = 32'd31856;
			33681: outdata = 32'd31855;
			33682: outdata = 32'd31854;
			33683: outdata = 32'd31853;
			33684: outdata = 32'd31852;
			33685: outdata = 32'd31851;
			33686: outdata = 32'd31850;
			33687: outdata = 32'd31849;
			33688: outdata = 32'd31848;
			33689: outdata = 32'd31847;
			33690: outdata = 32'd31846;
			33691: outdata = 32'd31845;
			33692: outdata = 32'd31844;
			33693: outdata = 32'd31843;
			33694: outdata = 32'd31842;
			33695: outdata = 32'd31841;
			33696: outdata = 32'd31840;
			33697: outdata = 32'd31839;
			33698: outdata = 32'd31838;
			33699: outdata = 32'd31837;
			33700: outdata = 32'd31836;
			33701: outdata = 32'd31835;
			33702: outdata = 32'd31834;
			33703: outdata = 32'd31833;
			33704: outdata = 32'd31832;
			33705: outdata = 32'd31831;
			33706: outdata = 32'd31830;
			33707: outdata = 32'd31829;
			33708: outdata = 32'd31828;
			33709: outdata = 32'd31827;
			33710: outdata = 32'd31826;
			33711: outdata = 32'd31825;
			33712: outdata = 32'd31824;
			33713: outdata = 32'd31823;
			33714: outdata = 32'd31822;
			33715: outdata = 32'd31821;
			33716: outdata = 32'd31820;
			33717: outdata = 32'd31819;
			33718: outdata = 32'd31818;
			33719: outdata = 32'd31817;
			33720: outdata = 32'd31816;
			33721: outdata = 32'd31815;
			33722: outdata = 32'd31814;
			33723: outdata = 32'd31813;
			33724: outdata = 32'd31812;
			33725: outdata = 32'd31811;
			33726: outdata = 32'd31810;
			33727: outdata = 32'd31809;
			33728: outdata = 32'd31808;
			33729: outdata = 32'd31807;
			33730: outdata = 32'd31806;
			33731: outdata = 32'd31805;
			33732: outdata = 32'd31804;
			33733: outdata = 32'd31803;
			33734: outdata = 32'd31802;
			33735: outdata = 32'd31801;
			33736: outdata = 32'd31800;
			33737: outdata = 32'd31799;
			33738: outdata = 32'd31798;
			33739: outdata = 32'd31797;
			33740: outdata = 32'd31796;
			33741: outdata = 32'd31795;
			33742: outdata = 32'd31794;
			33743: outdata = 32'd31793;
			33744: outdata = 32'd31792;
			33745: outdata = 32'd31791;
			33746: outdata = 32'd31790;
			33747: outdata = 32'd31789;
			33748: outdata = 32'd31788;
			33749: outdata = 32'd31787;
			33750: outdata = 32'd31786;
			33751: outdata = 32'd31785;
			33752: outdata = 32'd31784;
			33753: outdata = 32'd31783;
			33754: outdata = 32'd31782;
			33755: outdata = 32'd31781;
			33756: outdata = 32'd31780;
			33757: outdata = 32'd31779;
			33758: outdata = 32'd31778;
			33759: outdata = 32'd31777;
			33760: outdata = 32'd31776;
			33761: outdata = 32'd31775;
			33762: outdata = 32'd31774;
			33763: outdata = 32'd31773;
			33764: outdata = 32'd31772;
			33765: outdata = 32'd31771;
			33766: outdata = 32'd31770;
			33767: outdata = 32'd31769;
			33768: outdata = 32'd31768;
			33769: outdata = 32'd31767;
			33770: outdata = 32'd31766;
			33771: outdata = 32'd31765;
			33772: outdata = 32'd31764;
			33773: outdata = 32'd31763;
			33774: outdata = 32'd31762;
			33775: outdata = 32'd31761;
			33776: outdata = 32'd31760;
			33777: outdata = 32'd31759;
			33778: outdata = 32'd31758;
			33779: outdata = 32'd31757;
			33780: outdata = 32'd31756;
			33781: outdata = 32'd31755;
			33782: outdata = 32'd31754;
			33783: outdata = 32'd31753;
			33784: outdata = 32'd31752;
			33785: outdata = 32'd31751;
			33786: outdata = 32'd31750;
			33787: outdata = 32'd31749;
			33788: outdata = 32'd31748;
			33789: outdata = 32'd31747;
			33790: outdata = 32'd31746;
			33791: outdata = 32'd31745;
			33792: outdata = 32'd31744;
			33793: outdata = 32'd31743;
			33794: outdata = 32'd31742;
			33795: outdata = 32'd31741;
			33796: outdata = 32'd31740;
			33797: outdata = 32'd31739;
			33798: outdata = 32'd31738;
			33799: outdata = 32'd31737;
			33800: outdata = 32'd31736;
			33801: outdata = 32'd31735;
			33802: outdata = 32'd31734;
			33803: outdata = 32'd31733;
			33804: outdata = 32'd31732;
			33805: outdata = 32'd31731;
			33806: outdata = 32'd31730;
			33807: outdata = 32'd31729;
			33808: outdata = 32'd31728;
			33809: outdata = 32'd31727;
			33810: outdata = 32'd31726;
			33811: outdata = 32'd31725;
			33812: outdata = 32'd31724;
			33813: outdata = 32'd31723;
			33814: outdata = 32'd31722;
			33815: outdata = 32'd31721;
			33816: outdata = 32'd31720;
			33817: outdata = 32'd31719;
			33818: outdata = 32'd31718;
			33819: outdata = 32'd31717;
			33820: outdata = 32'd31716;
			33821: outdata = 32'd31715;
			33822: outdata = 32'd31714;
			33823: outdata = 32'd31713;
			33824: outdata = 32'd31712;
			33825: outdata = 32'd31711;
			33826: outdata = 32'd31710;
			33827: outdata = 32'd31709;
			33828: outdata = 32'd31708;
			33829: outdata = 32'd31707;
			33830: outdata = 32'd31706;
			33831: outdata = 32'd31705;
			33832: outdata = 32'd31704;
			33833: outdata = 32'd31703;
			33834: outdata = 32'd31702;
			33835: outdata = 32'd31701;
			33836: outdata = 32'd31700;
			33837: outdata = 32'd31699;
			33838: outdata = 32'd31698;
			33839: outdata = 32'd31697;
			33840: outdata = 32'd31696;
			33841: outdata = 32'd31695;
			33842: outdata = 32'd31694;
			33843: outdata = 32'd31693;
			33844: outdata = 32'd31692;
			33845: outdata = 32'd31691;
			33846: outdata = 32'd31690;
			33847: outdata = 32'd31689;
			33848: outdata = 32'd31688;
			33849: outdata = 32'd31687;
			33850: outdata = 32'd31686;
			33851: outdata = 32'd31685;
			33852: outdata = 32'd31684;
			33853: outdata = 32'd31683;
			33854: outdata = 32'd31682;
			33855: outdata = 32'd31681;
			33856: outdata = 32'd31680;
			33857: outdata = 32'd31679;
			33858: outdata = 32'd31678;
			33859: outdata = 32'd31677;
			33860: outdata = 32'd31676;
			33861: outdata = 32'd31675;
			33862: outdata = 32'd31674;
			33863: outdata = 32'd31673;
			33864: outdata = 32'd31672;
			33865: outdata = 32'd31671;
			33866: outdata = 32'd31670;
			33867: outdata = 32'd31669;
			33868: outdata = 32'd31668;
			33869: outdata = 32'd31667;
			33870: outdata = 32'd31666;
			33871: outdata = 32'd31665;
			33872: outdata = 32'd31664;
			33873: outdata = 32'd31663;
			33874: outdata = 32'd31662;
			33875: outdata = 32'd31661;
			33876: outdata = 32'd31660;
			33877: outdata = 32'd31659;
			33878: outdata = 32'd31658;
			33879: outdata = 32'd31657;
			33880: outdata = 32'd31656;
			33881: outdata = 32'd31655;
			33882: outdata = 32'd31654;
			33883: outdata = 32'd31653;
			33884: outdata = 32'd31652;
			33885: outdata = 32'd31651;
			33886: outdata = 32'd31650;
			33887: outdata = 32'd31649;
			33888: outdata = 32'd31648;
			33889: outdata = 32'd31647;
			33890: outdata = 32'd31646;
			33891: outdata = 32'd31645;
			33892: outdata = 32'd31644;
			33893: outdata = 32'd31643;
			33894: outdata = 32'd31642;
			33895: outdata = 32'd31641;
			33896: outdata = 32'd31640;
			33897: outdata = 32'd31639;
			33898: outdata = 32'd31638;
			33899: outdata = 32'd31637;
			33900: outdata = 32'd31636;
			33901: outdata = 32'd31635;
			33902: outdata = 32'd31634;
			33903: outdata = 32'd31633;
			33904: outdata = 32'd31632;
			33905: outdata = 32'd31631;
			33906: outdata = 32'd31630;
			33907: outdata = 32'd31629;
			33908: outdata = 32'd31628;
			33909: outdata = 32'd31627;
			33910: outdata = 32'd31626;
			33911: outdata = 32'd31625;
			33912: outdata = 32'd31624;
			33913: outdata = 32'd31623;
			33914: outdata = 32'd31622;
			33915: outdata = 32'd31621;
			33916: outdata = 32'd31620;
			33917: outdata = 32'd31619;
			33918: outdata = 32'd31618;
			33919: outdata = 32'd31617;
			33920: outdata = 32'd31616;
			33921: outdata = 32'd31615;
			33922: outdata = 32'd31614;
			33923: outdata = 32'd31613;
			33924: outdata = 32'd31612;
			33925: outdata = 32'd31611;
			33926: outdata = 32'd31610;
			33927: outdata = 32'd31609;
			33928: outdata = 32'd31608;
			33929: outdata = 32'd31607;
			33930: outdata = 32'd31606;
			33931: outdata = 32'd31605;
			33932: outdata = 32'd31604;
			33933: outdata = 32'd31603;
			33934: outdata = 32'd31602;
			33935: outdata = 32'd31601;
			33936: outdata = 32'd31600;
			33937: outdata = 32'd31599;
			33938: outdata = 32'd31598;
			33939: outdata = 32'd31597;
			33940: outdata = 32'd31596;
			33941: outdata = 32'd31595;
			33942: outdata = 32'd31594;
			33943: outdata = 32'd31593;
			33944: outdata = 32'd31592;
			33945: outdata = 32'd31591;
			33946: outdata = 32'd31590;
			33947: outdata = 32'd31589;
			33948: outdata = 32'd31588;
			33949: outdata = 32'd31587;
			33950: outdata = 32'd31586;
			33951: outdata = 32'd31585;
			33952: outdata = 32'd31584;
			33953: outdata = 32'd31583;
			33954: outdata = 32'd31582;
			33955: outdata = 32'd31581;
			33956: outdata = 32'd31580;
			33957: outdata = 32'd31579;
			33958: outdata = 32'd31578;
			33959: outdata = 32'd31577;
			33960: outdata = 32'd31576;
			33961: outdata = 32'd31575;
			33962: outdata = 32'd31574;
			33963: outdata = 32'd31573;
			33964: outdata = 32'd31572;
			33965: outdata = 32'd31571;
			33966: outdata = 32'd31570;
			33967: outdata = 32'd31569;
			33968: outdata = 32'd31568;
			33969: outdata = 32'd31567;
			33970: outdata = 32'd31566;
			33971: outdata = 32'd31565;
			33972: outdata = 32'd31564;
			33973: outdata = 32'd31563;
			33974: outdata = 32'd31562;
			33975: outdata = 32'd31561;
			33976: outdata = 32'd31560;
			33977: outdata = 32'd31559;
			33978: outdata = 32'd31558;
			33979: outdata = 32'd31557;
			33980: outdata = 32'd31556;
			33981: outdata = 32'd31555;
			33982: outdata = 32'd31554;
			33983: outdata = 32'd31553;
			33984: outdata = 32'd31552;
			33985: outdata = 32'd31551;
			33986: outdata = 32'd31550;
			33987: outdata = 32'd31549;
			33988: outdata = 32'd31548;
			33989: outdata = 32'd31547;
			33990: outdata = 32'd31546;
			33991: outdata = 32'd31545;
			33992: outdata = 32'd31544;
			33993: outdata = 32'd31543;
			33994: outdata = 32'd31542;
			33995: outdata = 32'd31541;
			33996: outdata = 32'd31540;
			33997: outdata = 32'd31539;
			33998: outdata = 32'd31538;
			33999: outdata = 32'd31537;
			34000: outdata = 32'd31536;
			34001: outdata = 32'd31535;
			34002: outdata = 32'd31534;
			34003: outdata = 32'd31533;
			34004: outdata = 32'd31532;
			34005: outdata = 32'd31531;
			34006: outdata = 32'd31530;
			34007: outdata = 32'd31529;
			34008: outdata = 32'd31528;
			34009: outdata = 32'd31527;
			34010: outdata = 32'd31526;
			34011: outdata = 32'd31525;
			34012: outdata = 32'd31524;
			34013: outdata = 32'd31523;
			34014: outdata = 32'd31522;
			34015: outdata = 32'd31521;
			34016: outdata = 32'd31520;
			34017: outdata = 32'd31519;
			34018: outdata = 32'd31518;
			34019: outdata = 32'd31517;
			34020: outdata = 32'd31516;
			34021: outdata = 32'd31515;
			34022: outdata = 32'd31514;
			34023: outdata = 32'd31513;
			34024: outdata = 32'd31512;
			34025: outdata = 32'd31511;
			34026: outdata = 32'd31510;
			34027: outdata = 32'd31509;
			34028: outdata = 32'd31508;
			34029: outdata = 32'd31507;
			34030: outdata = 32'd31506;
			34031: outdata = 32'd31505;
			34032: outdata = 32'd31504;
			34033: outdata = 32'd31503;
			34034: outdata = 32'd31502;
			34035: outdata = 32'd31501;
			34036: outdata = 32'd31500;
			34037: outdata = 32'd31499;
			34038: outdata = 32'd31498;
			34039: outdata = 32'd31497;
			34040: outdata = 32'd31496;
			34041: outdata = 32'd31495;
			34042: outdata = 32'd31494;
			34043: outdata = 32'd31493;
			34044: outdata = 32'd31492;
			34045: outdata = 32'd31491;
			34046: outdata = 32'd31490;
			34047: outdata = 32'd31489;
			34048: outdata = 32'd31488;
			34049: outdata = 32'd31487;
			34050: outdata = 32'd31486;
			34051: outdata = 32'd31485;
			34052: outdata = 32'd31484;
			34053: outdata = 32'd31483;
			34054: outdata = 32'd31482;
			34055: outdata = 32'd31481;
			34056: outdata = 32'd31480;
			34057: outdata = 32'd31479;
			34058: outdata = 32'd31478;
			34059: outdata = 32'd31477;
			34060: outdata = 32'd31476;
			34061: outdata = 32'd31475;
			34062: outdata = 32'd31474;
			34063: outdata = 32'd31473;
			34064: outdata = 32'd31472;
			34065: outdata = 32'd31471;
			34066: outdata = 32'd31470;
			34067: outdata = 32'd31469;
			34068: outdata = 32'd31468;
			34069: outdata = 32'd31467;
			34070: outdata = 32'd31466;
			34071: outdata = 32'd31465;
			34072: outdata = 32'd31464;
			34073: outdata = 32'd31463;
			34074: outdata = 32'd31462;
			34075: outdata = 32'd31461;
			34076: outdata = 32'd31460;
			34077: outdata = 32'd31459;
			34078: outdata = 32'd31458;
			34079: outdata = 32'd31457;
			34080: outdata = 32'd31456;
			34081: outdata = 32'd31455;
			34082: outdata = 32'd31454;
			34083: outdata = 32'd31453;
			34084: outdata = 32'd31452;
			34085: outdata = 32'd31451;
			34086: outdata = 32'd31450;
			34087: outdata = 32'd31449;
			34088: outdata = 32'd31448;
			34089: outdata = 32'd31447;
			34090: outdata = 32'd31446;
			34091: outdata = 32'd31445;
			34092: outdata = 32'd31444;
			34093: outdata = 32'd31443;
			34094: outdata = 32'd31442;
			34095: outdata = 32'd31441;
			34096: outdata = 32'd31440;
			34097: outdata = 32'd31439;
			34098: outdata = 32'd31438;
			34099: outdata = 32'd31437;
			34100: outdata = 32'd31436;
			34101: outdata = 32'd31435;
			34102: outdata = 32'd31434;
			34103: outdata = 32'd31433;
			34104: outdata = 32'd31432;
			34105: outdata = 32'd31431;
			34106: outdata = 32'd31430;
			34107: outdata = 32'd31429;
			34108: outdata = 32'd31428;
			34109: outdata = 32'd31427;
			34110: outdata = 32'd31426;
			34111: outdata = 32'd31425;
			34112: outdata = 32'd31424;
			34113: outdata = 32'd31423;
			34114: outdata = 32'd31422;
			34115: outdata = 32'd31421;
			34116: outdata = 32'd31420;
			34117: outdata = 32'd31419;
			34118: outdata = 32'd31418;
			34119: outdata = 32'd31417;
			34120: outdata = 32'd31416;
			34121: outdata = 32'd31415;
			34122: outdata = 32'd31414;
			34123: outdata = 32'd31413;
			34124: outdata = 32'd31412;
			34125: outdata = 32'd31411;
			34126: outdata = 32'd31410;
			34127: outdata = 32'd31409;
			34128: outdata = 32'd31408;
			34129: outdata = 32'd31407;
			34130: outdata = 32'd31406;
			34131: outdata = 32'd31405;
			34132: outdata = 32'd31404;
			34133: outdata = 32'd31403;
			34134: outdata = 32'd31402;
			34135: outdata = 32'd31401;
			34136: outdata = 32'd31400;
			34137: outdata = 32'd31399;
			34138: outdata = 32'd31398;
			34139: outdata = 32'd31397;
			34140: outdata = 32'd31396;
			34141: outdata = 32'd31395;
			34142: outdata = 32'd31394;
			34143: outdata = 32'd31393;
			34144: outdata = 32'd31392;
			34145: outdata = 32'd31391;
			34146: outdata = 32'd31390;
			34147: outdata = 32'd31389;
			34148: outdata = 32'd31388;
			34149: outdata = 32'd31387;
			34150: outdata = 32'd31386;
			34151: outdata = 32'd31385;
			34152: outdata = 32'd31384;
			34153: outdata = 32'd31383;
			34154: outdata = 32'd31382;
			34155: outdata = 32'd31381;
			34156: outdata = 32'd31380;
			34157: outdata = 32'd31379;
			34158: outdata = 32'd31378;
			34159: outdata = 32'd31377;
			34160: outdata = 32'd31376;
			34161: outdata = 32'd31375;
			34162: outdata = 32'd31374;
			34163: outdata = 32'd31373;
			34164: outdata = 32'd31372;
			34165: outdata = 32'd31371;
			34166: outdata = 32'd31370;
			34167: outdata = 32'd31369;
			34168: outdata = 32'd31368;
			34169: outdata = 32'd31367;
			34170: outdata = 32'd31366;
			34171: outdata = 32'd31365;
			34172: outdata = 32'd31364;
			34173: outdata = 32'd31363;
			34174: outdata = 32'd31362;
			34175: outdata = 32'd31361;
			34176: outdata = 32'd31360;
			34177: outdata = 32'd31359;
			34178: outdata = 32'd31358;
			34179: outdata = 32'd31357;
			34180: outdata = 32'd31356;
			34181: outdata = 32'd31355;
			34182: outdata = 32'd31354;
			34183: outdata = 32'd31353;
			34184: outdata = 32'd31352;
			34185: outdata = 32'd31351;
			34186: outdata = 32'd31350;
			34187: outdata = 32'd31349;
			34188: outdata = 32'd31348;
			34189: outdata = 32'd31347;
			34190: outdata = 32'd31346;
			34191: outdata = 32'd31345;
			34192: outdata = 32'd31344;
			34193: outdata = 32'd31343;
			34194: outdata = 32'd31342;
			34195: outdata = 32'd31341;
			34196: outdata = 32'd31340;
			34197: outdata = 32'd31339;
			34198: outdata = 32'd31338;
			34199: outdata = 32'd31337;
			34200: outdata = 32'd31336;
			34201: outdata = 32'd31335;
			34202: outdata = 32'd31334;
			34203: outdata = 32'd31333;
			34204: outdata = 32'd31332;
			34205: outdata = 32'd31331;
			34206: outdata = 32'd31330;
			34207: outdata = 32'd31329;
			34208: outdata = 32'd31328;
			34209: outdata = 32'd31327;
			34210: outdata = 32'd31326;
			34211: outdata = 32'd31325;
			34212: outdata = 32'd31324;
			34213: outdata = 32'd31323;
			34214: outdata = 32'd31322;
			34215: outdata = 32'd31321;
			34216: outdata = 32'd31320;
			34217: outdata = 32'd31319;
			34218: outdata = 32'd31318;
			34219: outdata = 32'd31317;
			34220: outdata = 32'd31316;
			34221: outdata = 32'd31315;
			34222: outdata = 32'd31314;
			34223: outdata = 32'd31313;
			34224: outdata = 32'd31312;
			34225: outdata = 32'd31311;
			34226: outdata = 32'd31310;
			34227: outdata = 32'd31309;
			34228: outdata = 32'd31308;
			34229: outdata = 32'd31307;
			34230: outdata = 32'd31306;
			34231: outdata = 32'd31305;
			34232: outdata = 32'd31304;
			34233: outdata = 32'd31303;
			34234: outdata = 32'd31302;
			34235: outdata = 32'd31301;
			34236: outdata = 32'd31300;
			34237: outdata = 32'd31299;
			34238: outdata = 32'd31298;
			34239: outdata = 32'd31297;
			34240: outdata = 32'd31296;
			34241: outdata = 32'd31295;
			34242: outdata = 32'd31294;
			34243: outdata = 32'd31293;
			34244: outdata = 32'd31292;
			34245: outdata = 32'd31291;
			34246: outdata = 32'd31290;
			34247: outdata = 32'd31289;
			34248: outdata = 32'd31288;
			34249: outdata = 32'd31287;
			34250: outdata = 32'd31286;
			34251: outdata = 32'd31285;
			34252: outdata = 32'd31284;
			34253: outdata = 32'd31283;
			34254: outdata = 32'd31282;
			34255: outdata = 32'd31281;
			34256: outdata = 32'd31280;
			34257: outdata = 32'd31279;
			34258: outdata = 32'd31278;
			34259: outdata = 32'd31277;
			34260: outdata = 32'd31276;
			34261: outdata = 32'd31275;
			34262: outdata = 32'd31274;
			34263: outdata = 32'd31273;
			34264: outdata = 32'd31272;
			34265: outdata = 32'd31271;
			34266: outdata = 32'd31270;
			34267: outdata = 32'd31269;
			34268: outdata = 32'd31268;
			34269: outdata = 32'd31267;
			34270: outdata = 32'd31266;
			34271: outdata = 32'd31265;
			34272: outdata = 32'd31264;
			34273: outdata = 32'd31263;
			34274: outdata = 32'd31262;
			34275: outdata = 32'd31261;
			34276: outdata = 32'd31260;
			34277: outdata = 32'd31259;
			34278: outdata = 32'd31258;
			34279: outdata = 32'd31257;
			34280: outdata = 32'd31256;
			34281: outdata = 32'd31255;
			34282: outdata = 32'd31254;
			34283: outdata = 32'd31253;
			34284: outdata = 32'd31252;
			34285: outdata = 32'd31251;
			34286: outdata = 32'd31250;
			34287: outdata = 32'd31249;
			34288: outdata = 32'd31248;
			34289: outdata = 32'd31247;
			34290: outdata = 32'd31246;
			34291: outdata = 32'd31245;
			34292: outdata = 32'd31244;
			34293: outdata = 32'd31243;
			34294: outdata = 32'd31242;
			34295: outdata = 32'd31241;
			34296: outdata = 32'd31240;
			34297: outdata = 32'd31239;
			34298: outdata = 32'd31238;
			34299: outdata = 32'd31237;
			34300: outdata = 32'd31236;
			34301: outdata = 32'd31235;
			34302: outdata = 32'd31234;
			34303: outdata = 32'd31233;
			34304: outdata = 32'd31232;
			34305: outdata = 32'd31231;
			34306: outdata = 32'd31230;
			34307: outdata = 32'd31229;
			34308: outdata = 32'd31228;
			34309: outdata = 32'd31227;
			34310: outdata = 32'd31226;
			34311: outdata = 32'd31225;
			34312: outdata = 32'd31224;
			34313: outdata = 32'd31223;
			34314: outdata = 32'd31222;
			34315: outdata = 32'd31221;
			34316: outdata = 32'd31220;
			34317: outdata = 32'd31219;
			34318: outdata = 32'd31218;
			34319: outdata = 32'd31217;
			34320: outdata = 32'd31216;
			34321: outdata = 32'd31215;
			34322: outdata = 32'd31214;
			34323: outdata = 32'd31213;
			34324: outdata = 32'd31212;
			34325: outdata = 32'd31211;
			34326: outdata = 32'd31210;
			34327: outdata = 32'd31209;
			34328: outdata = 32'd31208;
			34329: outdata = 32'd31207;
			34330: outdata = 32'd31206;
			34331: outdata = 32'd31205;
			34332: outdata = 32'd31204;
			34333: outdata = 32'd31203;
			34334: outdata = 32'd31202;
			34335: outdata = 32'd31201;
			34336: outdata = 32'd31200;
			34337: outdata = 32'd31199;
			34338: outdata = 32'd31198;
			34339: outdata = 32'd31197;
			34340: outdata = 32'd31196;
			34341: outdata = 32'd31195;
			34342: outdata = 32'd31194;
			34343: outdata = 32'd31193;
			34344: outdata = 32'd31192;
			34345: outdata = 32'd31191;
			34346: outdata = 32'd31190;
			34347: outdata = 32'd31189;
			34348: outdata = 32'd31188;
			34349: outdata = 32'd31187;
			34350: outdata = 32'd31186;
			34351: outdata = 32'd31185;
			34352: outdata = 32'd31184;
			34353: outdata = 32'd31183;
			34354: outdata = 32'd31182;
			34355: outdata = 32'd31181;
			34356: outdata = 32'd31180;
			34357: outdata = 32'd31179;
			34358: outdata = 32'd31178;
			34359: outdata = 32'd31177;
			34360: outdata = 32'd31176;
			34361: outdata = 32'd31175;
			34362: outdata = 32'd31174;
			34363: outdata = 32'd31173;
			34364: outdata = 32'd31172;
			34365: outdata = 32'd31171;
			34366: outdata = 32'd31170;
			34367: outdata = 32'd31169;
			34368: outdata = 32'd31168;
			34369: outdata = 32'd31167;
			34370: outdata = 32'd31166;
			34371: outdata = 32'd31165;
			34372: outdata = 32'd31164;
			34373: outdata = 32'd31163;
			34374: outdata = 32'd31162;
			34375: outdata = 32'd31161;
			34376: outdata = 32'd31160;
			34377: outdata = 32'd31159;
			34378: outdata = 32'd31158;
			34379: outdata = 32'd31157;
			34380: outdata = 32'd31156;
			34381: outdata = 32'd31155;
			34382: outdata = 32'd31154;
			34383: outdata = 32'd31153;
			34384: outdata = 32'd31152;
			34385: outdata = 32'd31151;
			34386: outdata = 32'd31150;
			34387: outdata = 32'd31149;
			34388: outdata = 32'd31148;
			34389: outdata = 32'd31147;
			34390: outdata = 32'd31146;
			34391: outdata = 32'd31145;
			34392: outdata = 32'd31144;
			34393: outdata = 32'd31143;
			34394: outdata = 32'd31142;
			34395: outdata = 32'd31141;
			34396: outdata = 32'd31140;
			34397: outdata = 32'd31139;
			34398: outdata = 32'd31138;
			34399: outdata = 32'd31137;
			34400: outdata = 32'd31136;
			34401: outdata = 32'd31135;
			34402: outdata = 32'd31134;
			34403: outdata = 32'd31133;
			34404: outdata = 32'd31132;
			34405: outdata = 32'd31131;
			34406: outdata = 32'd31130;
			34407: outdata = 32'd31129;
			34408: outdata = 32'd31128;
			34409: outdata = 32'd31127;
			34410: outdata = 32'd31126;
			34411: outdata = 32'd31125;
			34412: outdata = 32'd31124;
			34413: outdata = 32'd31123;
			34414: outdata = 32'd31122;
			34415: outdata = 32'd31121;
			34416: outdata = 32'd31120;
			34417: outdata = 32'd31119;
			34418: outdata = 32'd31118;
			34419: outdata = 32'd31117;
			34420: outdata = 32'd31116;
			34421: outdata = 32'd31115;
			34422: outdata = 32'd31114;
			34423: outdata = 32'd31113;
			34424: outdata = 32'd31112;
			34425: outdata = 32'd31111;
			34426: outdata = 32'd31110;
			34427: outdata = 32'd31109;
			34428: outdata = 32'd31108;
			34429: outdata = 32'd31107;
			34430: outdata = 32'd31106;
			34431: outdata = 32'd31105;
			34432: outdata = 32'd31104;
			34433: outdata = 32'd31103;
			34434: outdata = 32'd31102;
			34435: outdata = 32'd31101;
			34436: outdata = 32'd31100;
			34437: outdata = 32'd31099;
			34438: outdata = 32'd31098;
			34439: outdata = 32'd31097;
			34440: outdata = 32'd31096;
			34441: outdata = 32'd31095;
			34442: outdata = 32'd31094;
			34443: outdata = 32'd31093;
			34444: outdata = 32'd31092;
			34445: outdata = 32'd31091;
			34446: outdata = 32'd31090;
			34447: outdata = 32'd31089;
			34448: outdata = 32'd31088;
			34449: outdata = 32'd31087;
			34450: outdata = 32'd31086;
			34451: outdata = 32'd31085;
			34452: outdata = 32'd31084;
			34453: outdata = 32'd31083;
			34454: outdata = 32'd31082;
			34455: outdata = 32'd31081;
			34456: outdata = 32'd31080;
			34457: outdata = 32'd31079;
			34458: outdata = 32'd31078;
			34459: outdata = 32'd31077;
			34460: outdata = 32'd31076;
			34461: outdata = 32'd31075;
			34462: outdata = 32'd31074;
			34463: outdata = 32'd31073;
			34464: outdata = 32'd31072;
			34465: outdata = 32'd31071;
			34466: outdata = 32'd31070;
			34467: outdata = 32'd31069;
			34468: outdata = 32'd31068;
			34469: outdata = 32'd31067;
			34470: outdata = 32'd31066;
			34471: outdata = 32'd31065;
			34472: outdata = 32'd31064;
			34473: outdata = 32'd31063;
			34474: outdata = 32'd31062;
			34475: outdata = 32'd31061;
			34476: outdata = 32'd31060;
			34477: outdata = 32'd31059;
			34478: outdata = 32'd31058;
			34479: outdata = 32'd31057;
			34480: outdata = 32'd31056;
			34481: outdata = 32'd31055;
			34482: outdata = 32'd31054;
			34483: outdata = 32'd31053;
			34484: outdata = 32'd31052;
			34485: outdata = 32'd31051;
			34486: outdata = 32'd31050;
			34487: outdata = 32'd31049;
			34488: outdata = 32'd31048;
			34489: outdata = 32'd31047;
			34490: outdata = 32'd31046;
			34491: outdata = 32'd31045;
			34492: outdata = 32'd31044;
			34493: outdata = 32'd31043;
			34494: outdata = 32'd31042;
			34495: outdata = 32'd31041;
			34496: outdata = 32'd31040;
			34497: outdata = 32'd31039;
			34498: outdata = 32'd31038;
			34499: outdata = 32'd31037;
			34500: outdata = 32'd31036;
			34501: outdata = 32'd31035;
			34502: outdata = 32'd31034;
			34503: outdata = 32'd31033;
			34504: outdata = 32'd31032;
			34505: outdata = 32'd31031;
			34506: outdata = 32'd31030;
			34507: outdata = 32'd31029;
			34508: outdata = 32'd31028;
			34509: outdata = 32'd31027;
			34510: outdata = 32'd31026;
			34511: outdata = 32'd31025;
			34512: outdata = 32'd31024;
			34513: outdata = 32'd31023;
			34514: outdata = 32'd31022;
			34515: outdata = 32'd31021;
			34516: outdata = 32'd31020;
			34517: outdata = 32'd31019;
			34518: outdata = 32'd31018;
			34519: outdata = 32'd31017;
			34520: outdata = 32'd31016;
			34521: outdata = 32'd31015;
			34522: outdata = 32'd31014;
			34523: outdata = 32'd31013;
			34524: outdata = 32'd31012;
			34525: outdata = 32'd31011;
			34526: outdata = 32'd31010;
			34527: outdata = 32'd31009;
			34528: outdata = 32'd31008;
			34529: outdata = 32'd31007;
			34530: outdata = 32'd31006;
			34531: outdata = 32'd31005;
			34532: outdata = 32'd31004;
			34533: outdata = 32'd31003;
			34534: outdata = 32'd31002;
			34535: outdata = 32'd31001;
			34536: outdata = 32'd31000;
			34537: outdata = 32'd30999;
			34538: outdata = 32'd30998;
			34539: outdata = 32'd30997;
			34540: outdata = 32'd30996;
			34541: outdata = 32'd30995;
			34542: outdata = 32'd30994;
			34543: outdata = 32'd30993;
			34544: outdata = 32'd30992;
			34545: outdata = 32'd30991;
			34546: outdata = 32'd30990;
			34547: outdata = 32'd30989;
			34548: outdata = 32'd30988;
			34549: outdata = 32'd30987;
			34550: outdata = 32'd30986;
			34551: outdata = 32'd30985;
			34552: outdata = 32'd30984;
			34553: outdata = 32'd30983;
			34554: outdata = 32'd30982;
			34555: outdata = 32'd30981;
			34556: outdata = 32'd30980;
			34557: outdata = 32'd30979;
			34558: outdata = 32'd30978;
			34559: outdata = 32'd30977;
			34560: outdata = 32'd30976;
			34561: outdata = 32'd30975;
			34562: outdata = 32'd30974;
			34563: outdata = 32'd30973;
			34564: outdata = 32'd30972;
			34565: outdata = 32'd30971;
			34566: outdata = 32'd30970;
			34567: outdata = 32'd30969;
			34568: outdata = 32'd30968;
			34569: outdata = 32'd30967;
			34570: outdata = 32'd30966;
			34571: outdata = 32'd30965;
			34572: outdata = 32'd30964;
			34573: outdata = 32'd30963;
			34574: outdata = 32'd30962;
			34575: outdata = 32'd30961;
			34576: outdata = 32'd30960;
			34577: outdata = 32'd30959;
			34578: outdata = 32'd30958;
			34579: outdata = 32'd30957;
			34580: outdata = 32'd30956;
			34581: outdata = 32'd30955;
			34582: outdata = 32'd30954;
			34583: outdata = 32'd30953;
			34584: outdata = 32'd30952;
			34585: outdata = 32'd30951;
			34586: outdata = 32'd30950;
			34587: outdata = 32'd30949;
			34588: outdata = 32'd30948;
			34589: outdata = 32'd30947;
			34590: outdata = 32'd30946;
			34591: outdata = 32'd30945;
			34592: outdata = 32'd30944;
			34593: outdata = 32'd30943;
			34594: outdata = 32'd30942;
			34595: outdata = 32'd30941;
			34596: outdata = 32'd30940;
			34597: outdata = 32'd30939;
			34598: outdata = 32'd30938;
			34599: outdata = 32'd30937;
			34600: outdata = 32'd30936;
			34601: outdata = 32'd30935;
			34602: outdata = 32'd30934;
			34603: outdata = 32'd30933;
			34604: outdata = 32'd30932;
			34605: outdata = 32'd30931;
			34606: outdata = 32'd30930;
			34607: outdata = 32'd30929;
			34608: outdata = 32'd30928;
			34609: outdata = 32'd30927;
			34610: outdata = 32'd30926;
			34611: outdata = 32'd30925;
			34612: outdata = 32'd30924;
			34613: outdata = 32'd30923;
			34614: outdata = 32'd30922;
			34615: outdata = 32'd30921;
			34616: outdata = 32'd30920;
			34617: outdata = 32'd30919;
			34618: outdata = 32'd30918;
			34619: outdata = 32'd30917;
			34620: outdata = 32'd30916;
			34621: outdata = 32'd30915;
			34622: outdata = 32'd30914;
			34623: outdata = 32'd30913;
			34624: outdata = 32'd30912;
			34625: outdata = 32'd30911;
			34626: outdata = 32'd30910;
			34627: outdata = 32'd30909;
			34628: outdata = 32'd30908;
			34629: outdata = 32'd30907;
			34630: outdata = 32'd30906;
			34631: outdata = 32'd30905;
			34632: outdata = 32'd30904;
			34633: outdata = 32'd30903;
			34634: outdata = 32'd30902;
			34635: outdata = 32'd30901;
			34636: outdata = 32'd30900;
			34637: outdata = 32'd30899;
			34638: outdata = 32'd30898;
			34639: outdata = 32'd30897;
			34640: outdata = 32'd30896;
			34641: outdata = 32'd30895;
			34642: outdata = 32'd30894;
			34643: outdata = 32'd30893;
			34644: outdata = 32'd30892;
			34645: outdata = 32'd30891;
			34646: outdata = 32'd30890;
			34647: outdata = 32'd30889;
			34648: outdata = 32'd30888;
			34649: outdata = 32'd30887;
			34650: outdata = 32'd30886;
			34651: outdata = 32'd30885;
			34652: outdata = 32'd30884;
			34653: outdata = 32'd30883;
			34654: outdata = 32'd30882;
			34655: outdata = 32'd30881;
			34656: outdata = 32'd30880;
			34657: outdata = 32'd30879;
			34658: outdata = 32'd30878;
			34659: outdata = 32'd30877;
			34660: outdata = 32'd30876;
			34661: outdata = 32'd30875;
			34662: outdata = 32'd30874;
			34663: outdata = 32'd30873;
			34664: outdata = 32'd30872;
			34665: outdata = 32'd30871;
			34666: outdata = 32'd30870;
			34667: outdata = 32'd30869;
			34668: outdata = 32'd30868;
			34669: outdata = 32'd30867;
			34670: outdata = 32'd30866;
			34671: outdata = 32'd30865;
			34672: outdata = 32'd30864;
			34673: outdata = 32'd30863;
			34674: outdata = 32'd30862;
			34675: outdata = 32'd30861;
			34676: outdata = 32'd30860;
			34677: outdata = 32'd30859;
			34678: outdata = 32'd30858;
			34679: outdata = 32'd30857;
			34680: outdata = 32'd30856;
			34681: outdata = 32'd30855;
			34682: outdata = 32'd30854;
			34683: outdata = 32'd30853;
			34684: outdata = 32'd30852;
			34685: outdata = 32'd30851;
			34686: outdata = 32'd30850;
			34687: outdata = 32'd30849;
			34688: outdata = 32'd30848;
			34689: outdata = 32'd30847;
			34690: outdata = 32'd30846;
			34691: outdata = 32'd30845;
			34692: outdata = 32'd30844;
			34693: outdata = 32'd30843;
			34694: outdata = 32'd30842;
			34695: outdata = 32'd30841;
			34696: outdata = 32'd30840;
			34697: outdata = 32'd30839;
			34698: outdata = 32'd30838;
			34699: outdata = 32'd30837;
			34700: outdata = 32'd30836;
			34701: outdata = 32'd30835;
			34702: outdata = 32'd30834;
			34703: outdata = 32'd30833;
			34704: outdata = 32'd30832;
			34705: outdata = 32'd30831;
			34706: outdata = 32'd30830;
			34707: outdata = 32'd30829;
			34708: outdata = 32'd30828;
			34709: outdata = 32'd30827;
			34710: outdata = 32'd30826;
			34711: outdata = 32'd30825;
			34712: outdata = 32'd30824;
			34713: outdata = 32'd30823;
			34714: outdata = 32'd30822;
			34715: outdata = 32'd30821;
			34716: outdata = 32'd30820;
			34717: outdata = 32'd30819;
			34718: outdata = 32'd30818;
			34719: outdata = 32'd30817;
			34720: outdata = 32'd30816;
			34721: outdata = 32'd30815;
			34722: outdata = 32'd30814;
			34723: outdata = 32'd30813;
			34724: outdata = 32'd30812;
			34725: outdata = 32'd30811;
			34726: outdata = 32'd30810;
			34727: outdata = 32'd30809;
			34728: outdata = 32'd30808;
			34729: outdata = 32'd30807;
			34730: outdata = 32'd30806;
			34731: outdata = 32'd30805;
			34732: outdata = 32'd30804;
			34733: outdata = 32'd30803;
			34734: outdata = 32'd30802;
			34735: outdata = 32'd30801;
			34736: outdata = 32'd30800;
			34737: outdata = 32'd30799;
			34738: outdata = 32'd30798;
			34739: outdata = 32'd30797;
			34740: outdata = 32'd30796;
			34741: outdata = 32'd30795;
			34742: outdata = 32'd30794;
			34743: outdata = 32'd30793;
			34744: outdata = 32'd30792;
			34745: outdata = 32'd30791;
			34746: outdata = 32'd30790;
			34747: outdata = 32'd30789;
			34748: outdata = 32'd30788;
			34749: outdata = 32'd30787;
			34750: outdata = 32'd30786;
			34751: outdata = 32'd30785;
			34752: outdata = 32'd30784;
			34753: outdata = 32'd30783;
			34754: outdata = 32'd30782;
			34755: outdata = 32'd30781;
			34756: outdata = 32'd30780;
			34757: outdata = 32'd30779;
			34758: outdata = 32'd30778;
			34759: outdata = 32'd30777;
			34760: outdata = 32'd30776;
			34761: outdata = 32'd30775;
			34762: outdata = 32'd30774;
			34763: outdata = 32'd30773;
			34764: outdata = 32'd30772;
			34765: outdata = 32'd30771;
			34766: outdata = 32'd30770;
			34767: outdata = 32'd30769;
			34768: outdata = 32'd30768;
			34769: outdata = 32'd30767;
			34770: outdata = 32'd30766;
			34771: outdata = 32'd30765;
			34772: outdata = 32'd30764;
			34773: outdata = 32'd30763;
			34774: outdata = 32'd30762;
			34775: outdata = 32'd30761;
			34776: outdata = 32'd30760;
			34777: outdata = 32'd30759;
			34778: outdata = 32'd30758;
			34779: outdata = 32'd30757;
			34780: outdata = 32'd30756;
			34781: outdata = 32'd30755;
			34782: outdata = 32'd30754;
			34783: outdata = 32'd30753;
			34784: outdata = 32'd30752;
			34785: outdata = 32'd30751;
			34786: outdata = 32'd30750;
			34787: outdata = 32'd30749;
			34788: outdata = 32'd30748;
			34789: outdata = 32'd30747;
			34790: outdata = 32'd30746;
			34791: outdata = 32'd30745;
			34792: outdata = 32'd30744;
			34793: outdata = 32'd30743;
			34794: outdata = 32'd30742;
			34795: outdata = 32'd30741;
			34796: outdata = 32'd30740;
			34797: outdata = 32'd30739;
			34798: outdata = 32'd30738;
			34799: outdata = 32'd30737;
			34800: outdata = 32'd30736;
			34801: outdata = 32'd30735;
			34802: outdata = 32'd30734;
			34803: outdata = 32'd30733;
			34804: outdata = 32'd30732;
			34805: outdata = 32'd30731;
			34806: outdata = 32'd30730;
			34807: outdata = 32'd30729;
			34808: outdata = 32'd30728;
			34809: outdata = 32'd30727;
			34810: outdata = 32'd30726;
			34811: outdata = 32'd30725;
			34812: outdata = 32'd30724;
			34813: outdata = 32'd30723;
			34814: outdata = 32'd30722;
			34815: outdata = 32'd30721;
			34816: outdata = 32'd30720;
			34817: outdata = 32'd30719;
			34818: outdata = 32'd30718;
			34819: outdata = 32'd30717;
			34820: outdata = 32'd30716;
			34821: outdata = 32'd30715;
			34822: outdata = 32'd30714;
			34823: outdata = 32'd30713;
			34824: outdata = 32'd30712;
			34825: outdata = 32'd30711;
			34826: outdata = 32'd30710;
			34827: outdata = 32'd30709;
			34828: outdata = 32'd30708;
			34829: outdata = 32'd30707;
			34830: outdata = 32'd30706;
			34831: outdata = 32'd30705;
			34832: outdata = 32'd30704;
			34833: outdata = 32'd30703;
			34834: outdata = 32'd30702;
			34835: outdata = 32'd30701;
			34836: outdata = 32'd30700;
			34837: outdata = 32'd30699;
			34838: outdata = 32'd30698;
			34839: outdata = 32'd30697;
			34840: outdata = 32'd30696;
			34841: outdata = 32'd30695;
			34842: outdata = 32'd30694;
			34843: outdata = 32'd30693;
			34844: outdata = 32'd30692;
			34845: outdata = 32'd30691;
			34846: outdata = 32'd30690;
			34847: outdata = 32'd30689;
			34848: outdata = 32'd30688;
			34849: outdata = 32'd30687;
			34850: outdata = 32'd30686;
			34851: outdata = 32'd30685;
			34852: outdata = 32'd30684;
			34853: outdata = 32'd30683;
			34854: outdata = 32'd30682;
			34855: outdata = 32'd30681;
			34856: outdata = 32'd30680;
			34857: outdata = 32'd30679;
			34858: outdata = 32'd30678;
			34859: outdata = 32'd30677;
			34860: outdata = 32'd30676;
			34861: outdata = 32'd30675;
			34862: outdata = 32'd30674;
			34863: outdata = 32'd30673;
			34864: outdata = 32'd30672;
			34865: outdata = 32'd30671;
			34866: outdata = 32'd30670;
			34867: outdata = 32'd30669;
			34868: outdata = 32'd30668;
			34869: outdata = 32'd30667;
			34870: outdata = 32'd30666;
			34871: outdata = 32'd30665;
			34872: outdata = 32'd30664;
			34873: outdata = 32'd30663;
			34874: outdata = 32'd30662;
			34875: outdata = 32'd30661;
			34876: outdata = 32'd30660;
			34877: outdata = 32'd30659;
			34878: outdata = 32'd30658;
			34879: outdata = 32'd30657;
			34880: outdata = 32'd30656;
			34881: outdata = 32'd30655;
			34882: outdata = 32'd30654;
			34883: outdata = 32'd30653;
			34884: outdata = 32'd30652;
			34885: outdata = 32'd30651;
			34886: outdata = 32'd30650;
			34887: outdata = 32'd30649;
			34888: outdata = 32'd30648;
			34889: outdata = 32'd30647;
			34890: outdata = 32'd30646;
			34891: outdata = 32'd30645;
			34892: outdata = 32'd30644;
			34893: outdata = 32'd30643;
			34894: outdata = 32'd30642;
			34895: outdata = 32'd30641;
			34896: outdata = 32'd30640;
			34897: outdata = 32'd30639;
			34898: outdata = 32'd30638;
			34899: outdata = 32'd30637;
			34900: outdata = 32'd30636;
			34901: outdata = 32'd30635;
			34902: outdata = 32'd30634;
			34903: outdata = 32'd30633;
			34904: outdata = 32'd30632;
			34905: outdata = 32'd30631;
			34906: outdata = 32'd30630;
			34907: outdata = 32'd30629;
			34908: outdata = 32'd30628;
			34909: outdata = 32'd30627;
			34910: outdata = 32'd30626;
			34911: outdata = 32'd30625;
			34912: outdata = 32'd30624;
			34913: outdata = 32'd30623;
			34914: outdata = 32'd30622;
			34915: outdata = 32'd30621;
			34916: outdata = 32'd30620;
			34917: outdata = 32'd30619;
			34918: outdata = 32'd30618;
			34919: outdata = 32'd30617;
			34920: outdata = 32'd30616;
			34921: outdata = 32'd30615;
			34922: outdata = 32'd30614;
			34923: outdata = 32'd30613;
			34924: outdata = 32'd30612;
			34925: outdata = 32'd30611;
			34926: outdata = 32'd30610;
			34927: outdata = 32'd30609;
			34928: outdata = 32'd30608;
			34929: outdata = 32'd30607;
			34930: outdata = 32'd30606;
			34931: outdata = 32'd30605;
			34932: outdata = 32'd30604;
			34933: outdata = 32'd30603;
			34934: outdata = 32'd30602;
			34935: outdata = 32'd30601;
			34936: outdata = 32'd30600;
			34937: outdata = 32'd30599;
			34938: outdata = 32'd30598;
			34939: outdata = 32'd30597;
			34940: outdata = 32'd30596;
			34941: outdata = 32'd30595;
			34942: outdata = 32'd30594;
			34943: outdata = 32'd30593;
			34944: outdata = 32'd30592;
			34945: outdata = 32'd30591;
			34946: outdata = 32'd30590;
			34947: outdata = 32'd30589;
			34948: outdata = 32'd30588;
			34949: outdata = 32'd30587;
			34950: outdata = 32'd30586;
			34951: outdata = 32'd30585;
			34952: outdata = 32'd30584;
			34953: outdata = 32'd30583;
			34954: outdata = 32'd30582;
			34955: outdata = 32'd30581;
			34956: outdata = 32'd30580;
			34957: outdata = 32'd30579;
			34958: outdata = 32'd30578;
			34959: outdata = 32'd30577;
			34960: outdata = 32'd30576;
			34961: outdata = 32'd30575;
			34962: outdata = 32'd30574;
			34963: outdata = 32'd30573;
			34964: outdata = 32'd30572;
			34965: outdata = 32'd30571;
			34966: outdata = 32'd30570;
			34967: outdata = 32'd30569;
			34968: outdata = 32'd30568;
			34969: outdata = 32'd30567;
			34970: outdata = 32'd30566;
			34971: outdata = 32'd30565;
			34972: outdata = 32'd30564;
			34973: outdata = 32'd30563;
			34974: outdata = 32'd30562;
			34975: outdata = 32'd30561;
			34976: outdata = 32'd30560;
			34977: outdata = 32'd30559;
			34978: outdata = 32'd30558;
			34979: outdata = 32'd30557;
			34980: outdata = 32'd30556;
			34981: outdata = 32'd30555;
			34982: outdata = 32'd30554;
			34983: outdata = 32'd30553;
			34984: outdata = 32'd30552;
			34985: outdata = 32'd30551;
			34986: outdata = 32'd30550;
			34987: outdata = 32'd30549;
			34988: outdata = 32'd30548;
			34989: outdata = 32'd30547;
			34990: outdata = 32'd30546;
			34991: outdata = 32'd30545;
			34992: outdata = 32'd30544;
			34993: outdata = 32'd30543;
			34994: outdata = 32'd30542;
			34995: outdata = 32'd30541;
			34996: outdata = 32'd30540;
			34997: outdata = 32'd30539;
			34998: outdata = 32'd30538;
			34999: outdata = 32'd30537;
			35000: outdata = 32'd30536;
			35001: outdata = 32'd30535;
			35002: outdata = 32'd30534;
			35003: outdata = 32'd30533;
			35004: outdata = 32'd30532;
			35005: outdata = 32'd30531;
			35006: outdata = 32'd30530;
			35007: outdata = 32'd30529;
			35008: outdata = 32'd30528;
			35009: outdata = 32'd30527;
			35010: outdata = 32'd30526;
			35011: outdata = 32'd30525;
			35012: outdata = 32'd30524;
			35013: outdata = 32'd30523;
			35014: outdata = 32'd30522;
			35015: outdata = 32'd30521;
			35016: outdata = 32'd30520;
			35017: outdata = 32'd30519;
			35018: outdata = 32'd30518;
			35019: outdata = 32'd30517;
			35020: outdata = 32'd30516;
			35021: outdata = 32'd30515;
			35022: outdata = 32'd30514;
			35023: outdata = 32'd30513;
			35024: outdata = 32'd30512;
			35025: outdata = 32'd30511;
			35026: outdata = 32'd30510;
			35027: outdata = 32'd30509;
			35028: outdata = 32'd30508;
			35029: outdata = 32'd30507;
			35030: outdata = 32'd30506;
			35031: outdata = 32'd30505;
			35032: outdata = 32'd30504;
			35033: outdata = 32'd30503;
			35034: outdata = 32'd30502;
			35035: outdata = 32'd30501;
			35036: outdata = 32'd30500;
			35037: outdata = 32'd30499;
			35038: outdata = 32'd30498;
			35039: outdata = 32'd30497;
			35040: outdata = 32'd30496;
			35041: outdata = 32'd30495;
			35042: outdata = 32'd30494;
			35043: outdata = 32'd30493;
			35044: outdata = 32'd30492;
			35045: outdata = 32'd30491;
			35046: outdata = 32'd30490;
			35047: outdata = 32'd30489;
			35048: outdata = 32'd30488;
			35049: outdata = 32'd30487;
			35050: outdata = 32'd30486;
			35051: outdata = 32'd30485;
			35052: outdata = 32'd30484;
			35053: outdata = 32'd30483;
			35054: outdata = 32'd30482;
			35055: outdata = 32'd30481;
			35056: outdata = 32'd30480;
			35057: outdata = 32'd30479;
			35058: outdata = 32'd30478;
			35059: outdata = 32'd30477;
			35060: outdata = 32'd30476;
			35061: outdata = 32'd30475;
			35062: outdata = 32'd30474;
			35063: outdata = 32'd30473;
			35064: outdata = 32'd30472;
			35065: outdata = 32'd30471;
			35066: outdata = 32'd30470;
			35067: outdata = 32'd30469;
			35068: outdata = 32'd30468;
			35069: outdata = 32'd30467;
			35070: outdata = 32'd30466;
			35071: outdata = 32'd30465;
			35072: outdata = 32'd30464;
			35073: outdata = 32'd30463;
			35074: outdata = 32'd30462;
			35075: outdata = 32'd30461;
			35076: outdata = 32'd30460;
			35077: outdata = 32'd30459;
			35078: outdata = 32'd30458;
			35079: outdata = 32'd30457;
			35080: outdata = 32'd30456;
			35081: outdata = 32'd30455;
			35082: outdata = 32'd30454;
			35083: outdata = 32'd30453;
			35084: outdata = 32'd30452;
			35085: outdata = 32'd30451;
			35086: outdata = 32'd30450;
			35087: outdata = 32'd30449;
			35088: outdata = 32'd30448;
			35089: outdata = 32'd30447;
			35090: outdata = 32'd30446;
			35091: outdata = 32'd30445;
			35092: outdata = 32'd30444;
			35093: outdata = 32'd30443;
			35094: outdata = 32'd30442;
			35095: outdata = 32'd30441;
			35096: outdata = 32'd30440;
			35097: outdata = 32'd30439;
			35098: outdata = 32'd30438;
			35099: outdata = 32'd30437;
			35100: outdata = 32'd30436;
			35101: outdata = 32'd30435;
			35102: outdata = 32'd30434;
			35103: outdata = 32'd30433;
			35104: outdata = 32'd30432;
			35105: outdata = 32'd30431;
			35106: outdata = 32'd30430;
			35107: outdata = 32'd30429;
			35108: outdata = 32'd30428;
			35109: outdata = 32'd30427;
			35110: outdata = 32'd30426;
			35111: outdata = 32'd30425;
			35112: outdata = 32'd30424;
			35113: outdata = 32'd30423;
			35114: outdata = 32'd30422;
			35115: outdata = 32'd30421;
			35116: outdata = 32'd30420;
			35117: outdata = 32'd30419;
			35118: outdata = 32'd30418;
			35119: outdata = 32'd30417;
			35120: outdata = 32'd30416;
			35121: outdata = 32'd30415;
			35122: outdata = 32'd30414;
			35123: outdata = 32'd30413;
			35124: outdata = 32'd30412;
			35125: outdata = 32'd30411;
			35126: outdata = 32'd30410;
			35127: outdata = 32'd30409;
			35128: outdata = 32'd30408;
			35129: outdata = 32'd30407;
			35130: outdata = 32'd30406;
			35131: outdata = 32'd30405;
			35132: outdata = 32'd30404;
			35133: outdata = 32'd30403;
			35134: outdata = 32'd30402;
			35135: outdata = 32'd30401;
			35136: outdata = 32'd30400;
			35137: outdata = 32'd30399;
			35138: outdata = 32'd30398;
			35139: outdata = 32'd30397;
			35140: outdata = 32'd30396;
			35141: outdata = 32'd30395;
			35142: outdata = 32'd30394;
			35143: outdata = 32'd30393;
			35144: outdata = 32'd30392;
			35145: outdata = 32'd30391;
			35146: outdata = 32'd30390;
			35147: outdata = 32'd30389;
			35148: outdata = 32'd30388;
			35149: outdata = 32'd30387;
			35150: outdata = 32'd30386;
			35151: outdata = 32'd30385;
			35152: outdata = 32'd30384;
			35153: outdata = 32'd30383;
			35154: outdata = 32'd30382;
			35155: outdata = 32'd30381;
			35156: outdata = 32'd30380;
			35157: outdata = 32'd30379;
			35158: outdata = 32'd30378;
			35159: outdata = 32'd30377;
			35160: outdata = 32'd30376;
			35161: outdata = 32'd30375;
			35162: outdata = 32'd30374;
			35163: outdata = 32'd30373;
			35164: outdata = 32'd30372;
			35165: outdata = 32'd30371;
			35166: outdata = 32'd30370;
			35167: outdata = 32'd30369;
			35168: outdata = 32'd30368;
			35169: outdata = 32'd30367;
			35170: outdata = 32'd30366;
			35171: outdata = 32'd30365;
			35172: outdata = 32'd30364;
			35173: outdata = 32'd30363;
			35174: outdata = 32'd30362;
			35175: outdata = 32'd30361;
			35176: outdata = 32'd30360;
			35177: outdata = 32'd30359;
			35178: outdata = 32'd30358;
			35179: outdata = 32'd30357;
			35180: outdata = 32'd30356;
			35181: outdata = 32'd30355;
			35182: outdata = 32'd30354;
			35183: outdata = 32'd30353;
			35184: outdata = 32'd30352;
			35185: outdata = 32'd30351;
			35186: outdata = 32'd30350;
			35187: outdata = 32'd30349;
			35188: outdata = 32'd30348;
			35189: outdata = 32'd30347;
			35190: outdata = 32'd30346;
			35191: outdata = 32'd30345;
			35192: outdata = 32'd30344;
			35193: outdata = 32'd30343;
			35194: outdata = 32'd30342;
			35195: outdata = 32'd30341;
			35196: outdata = 32'd30340;
			35197: outdata = 32'd30339;
			35198: outdata = 32'd30338;
			35199: outdata = 32'd30337;
			35200: outdata = 32'd30336;
			35201: outdata = 32'd30335;
			35202: outdata = 32'd30334;
			35203: outdata = 32'd30333;
			35204: outdata = 32'd30332;
			35205: outdata = 32'd30331;
			35206: outdata = 32'd30330;
			35207: outdata = 32'd30329;
			35208: outdata = 32'd30328;
			35209: outdata = 32'd30327;
			35210: outdata = 32'd30326;
			35211: outdata = 32'd30325;
			35212: outdata = 32'd30324;
			35213: outdata = 32'd30323;
			35214: outdata = 32'd30322;
			35215: outdata = 32'd30321;
			35216: outdata = 32'd30320;
			35217: outdata = 32'd30319;
			35218: outdata = 32'd30318;
			35219: outdata = 32'd30317;
			35220: outdata = 32'd30316;
			35221: outdata = 32'd30315;
			35222: outdata = 32'd30314;
			35223: outdata = 32'd30313;
			35224: outdata = 32'd30312;
			35225: outdata = 32'd30311;
			35226: outdata = 32'd30310;
			35227: outdata = 32'd30309;
			35228: outdata = 32'd30308;
			35229: outdata = 32'd30307;
			35230: outdata = 32'd30306;
			35231: outdata = 32'd30305;
			35232: outdata = 32'd30304;
			35233: outdata = 32'd30303;
			35234: outdata = 32'd30302;
			35235: outdata = 32'd30301;
			35236: outdata = 32'd30300;
			35237: outdata = 32'd30299;
			35238: outdata = 32'd30298;
			35239: outdata = 32'd30297;
			35240: outdata = 32'd30296;
			35241: outdata = 32'd30295;
			35242: outdata = 32'd30294;
			35243: outdata = 32'd30293;
			35244: outdata = 32'd30292;
			35245: outdata = 32'd30291;
			35246: outdata = 32'd30290;
			35247: outdata = 32'd30289;
			35248: outdata = 32'd30288;
			35249: outdata = 32'd30287;
			35250: outdata = 32'd30286;
			35251: outdata = 32'd30285;
			35252: outdata = 32'd30284;
			35253: outdata = 32'd30283;
			35254: outdata = 32'd30282;
			35255: outdata = 32'd30281;
			35256: outdata = 32'd30280;
			35257: outdata = 32'd30279;
			35258: outdata = 32'd30278;
			35259: outdata = 32'd30277;
			35260: outdata = 32'd30276;
			35261: outdata = 32'd30275;
			35262: outdata = 32'd30274;
			35263: outdata = 32'd30273;
			35264: outdata = 32'd30272;
			35265: outdata = 32'd30271;
			35266: outdata = 32'd30270;
			35267: outdata = 32'd30269;
			35268: outdata = 32'd30268;
			35269: outdata = 32'd30267;
			35270: outdata = 32'd30266;
			35271: outdata = 32'd30265;
			35272: outdata = 32'd30264;
			35273: outdata = 32'd30263;
			35274: outdata = 32'd30262;
			35275: outdata = 32'd30261;
			35276: outdata = 32'd30260;
			35277: outdata = 32'd30259;
			35278: outdata = 32'd30258;
			35279: outdata = 32'd30257;
			35280: outdata = 32'd30256;
			35281: outdata = 32'd30255;
			35282: outdata = 32'd30254;
			35283: outdata = 32'd30253;
			35284: outdata = 32'd30252;
			35285: outdata = 32'd30251;
			35286: outdata = 32'd30250;
			35287: outdata = 32'd30249;
			35288: outdata = 32'd30248;
			35289: outdata = 32'd30247;
			35290: outdata = 32'd30246;
			35291: outdata = 32'd30245;
			35292: outdata = 32'd30244;
			35293: outdata = 32'd30243;
			35294: outdata = 32'd30242;
			35295: outdata = 32'd30241;
			35296: outdata = 32'd30240;
			35297: outdata = 32'd30239;
			35298: outdata = 32'd30238;
			35299: outdata = 32'd30237;
			35300: outdata = 32'd30236;
			35301: outdata = 32'd30235;
			35302: outdata = 32'd30234;
			35303: outdata = 32'd30233;
			35304: outdata = 32'd30232;
			35305: outdata = 32'd30231;
			35306: outdata = 32'd30230;
			35307: outdata = 32'd30229;
			35308: outdata = 32'd30228;
			35309: outdata = 32'd30227;
			35310: outdata = 32'd30226;
			35311: outdata = 32'd30225;
			35312: outdata = 32'd30224;
			35313: outdata = 32'd30223;
			35314: outdata = 32'd30222;
			35315: outdata = 32'd30221;
			35316: outdata = 32'd30220;
			35317: outdata = 32'd30219;
			35318: outdata = 32'd30218;
			35319: outdata = 32'd30217;
			35320: outdata = 32'd30216;
			35321: outdata = 32'd30215;
			35322: outdata = 32'd30214;
			35323: outdata = 32'd30213;
			35324: outdata = 32'd30212;
			35325: outdata = 32'd30211;
			35326: outdata = 32'd30210;
			35327: outdata = 32'd30209;
			35328: outdata = 32'd30208;
			35329: outdata = 32'd30207;
			35330: outdata = 32'd30206;
			35331: outdata = 32'd30205;
			35332: outdata = 32'd30204;
			35333: outdata = 32'd30203;
			35334: outdata = 32'd30202;
			35335: outdata = 32'd30201;
			35336: outdata = 32'd30200;
			35337: outdata = 32'd30199;
			35338: outdata = 32'd30198;
			35339: outdata = 32'd30197;
			35340: outdata = 32'd30196;
			35341: outdata = 32'd30195;
			35342: outdata = 32'd30194;
			35343: outdata = 32'd30193;
			35344: outdata = 32'd30192;
			35345: outdata = 32'd30191;
			35346: outdata = 32'd30190;
			35347: outdata = 32'd30189;
			35348: outdata = 32'd30188;
			35349: outdata = 32'd30187;
			35350: outdata = 32'd30186;
			35351: outdata = 32'd30185;
			35352: outdata = 32'd30184;
			35353: outdata = 32'd30183;
			35354: outdata = 32'd30182;
			35355: outdata = 32'd30181;
			35356: outdata = 32'd30180;
			35357: outdata = 32'd30179;
			35358: outdata = 32'd30178;
			35359: outdata = 32'd30177;
			35360: outdata = 32'd30176;
			35361: outdata = 32'd30175;
			35362: outdata = 32'd30174;
			35363: outdata = 32'd30173;
			35364: outdata = 32'd30172;
			35365: outdata = 32'd30171;
			35366: outdata = 32'd30170;
			35367: outdata = 32'd30169;
			35368: outdata = 32'd30168;
			35369: outdata = 32'd30167;
			35370: outdata = 32'd30166;
			35371: outdata = 32'd30165;
			35372: outdata = 32'd30164;
			35373: outdata = 32'd30163;
			35374: outdata = 32'd30162;
			35375: outdata = 32'd30161;
			35376: outdata = 32'd30160;
			35377: outdata = 32'd30159;
			35378: outdata = 32'd30158;
			35379: outdata = 32'd30157;
			35380: outdata = 32'd30156;
			35381: outdata = 32'd30155;
			35382: outdata = 32'd30154;
			35383: outdata = 32'd30153;
			35384: outdata = 32'd30152;
			35385: outdata = 32'd30151;
			35386: outdata = 32'd30150;
			35387: outdata = 32'd30149;
			35388: outdata = 32'd30148;
			35389: outdata = 32'd30147;
			35390: outdata = 32'd30146;
			35391: outdata = 32'd30145;
			35392: outdata = 32'd30144;
			35393: outdata = 32'd30143;
			35394: outdata = 32'd30142;
			35395: outdata = 32'd30141;
			35396: outdata = 32'd30140;
			35397: outdata = 32'd30139;
			35398: outdata = 32'd30138;
			35399: outdata = 32'd30137;
			35400: outdata = 32'd30136;
			35401: outdata = 32'd30135;
			35402: outdata = 32'd30134;
			35403: outdata = 32'd30133;
			35404: outdata = 32'd30132;
			35405: outdata = 32'd30131;
			35406: outdata = 32'd30130;
			35407: outdata = 32'd30129;
			35408: outdata = 32'd30128;
			35409: outdata = 32'd30127;
			35410: outdata = 32'd30126;
			35411: outdata = 32'd30125;
			35412: outdata = 32'd30124;
			35413: outdata = 32'd30123;
			35414: outdata = 32'd30122;
			35415: outdata = 32'd30121;
			35416: outdata = 32'd30120;
			35417: outdata = 32'd30119;
			35418: outdata = 32'd30118;
			35419: outdata = 32'd30117;
			35420: outdata = 32'd30116;
			35421: outdata = 32'd30115;
			35422: outdata = 32'd30114;
			35423: outdata = 32'd30113;
			35424: outdata = 32'd30112;
			35425: outdata = 32'd30111;
			35426: outdata = 32'd30110;
			35427: outdata = 32'd30109;
			35428: outdata = 32'd30108;
			35429: outdata = 32'd30107;
			35430: outdata = 32'd30106;
			35431: outdata = 32'd30105;
			35432: outdata = 32'd30104;
			35433: outdata = 32'd30103;
			35434: outdata = 32'd30102;
			35435: outdata = 32'd30101;
			35436: outdata = 32'd30100;
			35437: outdata = 32'd30099;
			35438: outdata = 32'd30098;
			35439: outdata = 32'd30097;
			35440: outdata = 32'd30096;
			35441: outdata = 32'd30095;
			35442: outdata = 32'd30094;
			35443: outdata = 32'd30093;
			35444: outdata = 32'd30092;
			35445: outdata = 32'd30091;
			35446: outdata = 32'd30090;
			35447: outdata = 32'd30089;
			35448: outdata = 32'd30088;
			35449: outdata = 32'd30087;
			35450: outdata = 32'd30086;
			35451: outdata = 32'd30085;
			35452: outdata = 32'd30084;
			35453: outdata = 32'd30083;
			35454: outdata = 32'd30082;
			35455: outdata = 32'd30081;
			35456: outdata = 32'd30080;
			35457: outdata = 32'd30079;
			35458: outdata = 32'd30078;
			35459: outdata = 32'd30077;
			35460: outdata = 32'd30076;
			35461: outdata = 32'd30075;
			35462: outdata = 32'd30074;
			35463: outdata = 32'd30073;
			35464: outdata = 32'd30072;
			35465: outdata = 32'd30071;
			35466: outdata = 32'd30070;
			35467: outdata = 32'd30069;
			35468: outdata = 32'd30068;
			35469: outdata = 32'd30067;
			35470: outdata = 32'd30066;
			35471: outdata = 32'd30065;
			35472: outdata = 32'd30064;
			35473: outdata = 32'd30063;
			35474: outdata = 32'd30062;
			35475: outdata = 32'd30061;
			35476: outdata = 32'd30060;
			35477: outdata = 32'd30059;
			35478: outdata = 32'd30058;
			35479: outdata = 32'd30057;
			35480: outdata = 32'd30056;
			35481: outdata = 32'd30055;
			35482: outdata = 32'd30054;
			35483: outdata = 32'd30053;
			35484: outdata = 32'd30052;
			35485: outdata = 32'd30051;
			35486: outdata = 32'd30050;
			35487: outdata = 32'd30049;
			35488: outdata = 32'd30048;
			35489: outdata = 32'd30047;
			35490: outdata = 32'd30046;
			35491: outdata = 32'd30045;
			35492: outdata = 32'd30044;
			35493: outdata = 32'd30043;
			35494: outdata = 32'd30042;
			35495: outdata = 32'd30041;
			35496: outdata = 32'd30040;
			35497: outdata = 32'd30039;
			35498: outdata = 32'd30038;
			35499: outdata = 32'd30037;
			35500: outdata = 32'd30036;
			35501: outdata = 32'd30035;
			35502: outdata = 32'd30034;
			35503: outdata = 32'd30033;
			35504: outdata = 32'd30032;
			35505: outdata = 32'd30031;
			35506: outdata = 32'd30030;
			35507: outdata = 32'd30029;
			35508: outdata = 32'd30028;
			35509: outdata = 32'd30027;
			35510: outdata = 32'd30026;
			35511: outdata = 32'd30025;
			35512: outdata = 32'd30024;
			35513: outdata = 32'd30023;
			35514: outdata = 32'd30022;
			35515: outdata = 32'd30021;
			35516: outdata = 32'd30020;
			35517: outdata = 32'd30019;
			35518: outdata = 32'd30018;
			35519: outdata = 32'd30017;
			35520: outdata = 32'd30016;
			35521: outdata = 32'd30015;
			35522: outdata = 32'd30014;
			35523: outdata = 32'd30013;
			35524: outdata = 32'd30012;
			35525: outdata = 32'd30011;
			35526: outdata = 32'd30010;
			35527: outdata = 32'd30009;
			35528: outdata = 32'd30008;
			35529: outdata = 32'd30007;
			35530: outdata = 32'd30006;
			35531: outdata = 32'd30005;
			35532: outdata = 32'd30004;
			35533: outdata = 32'd30003;
			35534: outdata = 32'd30002;
			35535: outdata = 32'd30001;
			35536: outdata = 32'd30000;
			35537: outdata = 32'd29999;
			35538: outdata = 32'd29998;
			35539: outdata = 32'd29997;
			35540: outdata = 32'd29996;
			35541: outdata = 32'd29995;
			35542: outdata = 32'd29994;
			35543: outdata = 32'd29993;
			35544: outdata = 32'd29992;
			35545: outdata = 32'd29991;
			35546: outdata = 32'd29990;
			35547: outdata = 32'd29989;
			35548: outdata = 32'd29988;
			35549: outdata = 32'd29987;
			35550: outdata = 32'd29986;
			35551: outdata = 32'd29985;
			35552: outdata = 32'd29984;
			35553: outdata = 32'd29983;
			35554: outdata = 32'd29982;
			35555: outdata = 32'd29981;
			35556: outdata = 32'd29980;
			35557: outdata = 32'd29979;
			35558: outdata = 32'd29978;
			35559: outdata = 32'd29977;
			35560: outdata = 32'd29976;
			35561: outdata = 32'd29975;
			35562: outdata = 32'd29974;
			35563: outdata = 32'd29973;
			35564: outdata = 32'd29972;
			35565: outdata = 32'd29971;
			35566: outdata = 32'd29970;
			35567: outdata = 32'd29969;
			35568: outdata = 32'd29968;
			35569: outdata = 32'd29967;
			35570: outdata = 32'd29966;
			35571: outdata = 32'd29965;
			35572: outdata = 32'd29964;
			35573: outdata = 32'd29963;
			35574: outdata = 32'd29962;
			35575: outdata = 32'd29961;
			35576: outdata = 32'd29960;
			35577: outdata = 32'd29959;
			35578: outdata = 32'd29958;
			35579: outdata = 32'd29957;
			35580: outdata = 32'd29956;
			35581: outdata = 32'd29955;
			35582: outdata = 32'd29954;
			35583: outdata = 32'd29953;
			35584: outdata = 32'd29952;
			35585: outdata = 32'd29951;
			35586: outdata = 32'd29950;
			35587: outdata = 32'd29949;
			35588: outdata = 32'd29948;
			35589: outdata = 32'd29947;
			35590: outdata = 32'd29946;
			35591: outdata = 32'd29945;
			35592: outdata = 32'd29944;
			35593: outdata = 32'd29943;
			35594: outdata = 32'd29942;
			35595: outdata = 32'd29941;
			35596: outdata = 32'd29940;
			35597: outdata = 32'd29939;
			35598: outdata = 32'd29938;
			35599: outdata = 32'd29937;
			35600: outdata = 32'd29936;
			35601: outdata = 32'd29935;
			35602: outdata = 32'd29934;
			35603: outdata = 32'd29933;
			35604: outdata = 32'd29932;
			35605: outdata = 32'd29931;
			35606: outdata = 32'd29930;
			35607: outdata = 32'd29929;
			35608: outdata = 32'd29928;
			35609: outdata = 32'd29927;
			35610: outdata = 32'd29926;
			35611: outdata = 32'd29925;
			35612: outdata = 32'd29924;
			35613: outdata = 32'd29923;
			35614: outdata = 32'd29922;
			35615: outdata = 32'd29921;
			35616: outdata = 32'd29920;
			35617: outdata = 32'd29919;
			35618: outdata = 32'd29918;
			35619: outdata = 32'd29917;
			35620: outdata = 32'd29916;
			35621: outdata = 32'd29915;
			35622: outdata = 32'd29914;
			35623: outdata = 32'd29913;
			35624: outdata = 32'd29912;
			35625: outdata = 32'd29911;
			35626: outdata = 32'd29910;
			35627: outdata = 32'd29909;
			35628: outdata = 32'd29908;
			35629: outdata = 32'd29907;
			35630: outdata = 32'd29906;
			35631: outdata = 32'd29905;
			35632: outdata = 32'd29904;
			35633: outdata = 32'd29903;
			35634: outdata = 32'd29902;
			35635: outdata = 32'd29901;
			35636: outdata = 32'd29900;
			35637: outdata = 32'd29899;
			35638: outdata = 32'd29898;
			35639: outdata = 32'd29897;
			35640: outdata = 32'd29896;
			35641: outdata = 32'd29895;
			35642: outdata = 32'd29894;
			35643: outdata = 32'd29893;
			35644: outdata = 32'd29892;
			35645: outdata = 32'd29891;
			35646: outdata = 32'd29890;
			35647: outdata = 32'd29889;
			35648: outdata = 32'd29888;
			35649: outdata = 32'd29887;
			35650: outdata = 32'd29886;
			35651: outdata = 32'd29885;
			35652: outdata = 32'd29884;
			35653: outdata = 32'd29883;
			35654: outdata = 32'd29882;
			35655: outdata = 32'd29881;
			35656: outdata = 32'd29880;
			35657: outdata = 32'd29879;
			35658: outdata = 32'd29878;
			35659: outdata = 32'd29877;
			35660: outdata = 32'd29876;
			35661: outdata = 32'd29875;
			35662: outdata = 32'd29874;
			35663: outdata = 32'd29873;
			35664: outdata = 32'd29872;
			35665: outdata = 32'd29871;
			35666: outdata = 32'd29870;
			35667: outdata = 32'd29869;
			35668: outdata = 32'd29868;
			35669: outdata = 32'd29867;
			35670: outdata = 32'd29866;
			35671: outdata = 32'd29865;
			35672: outdata = 32'd29864;
			35673: outdata = 32'd29863;
			35674: outdata = 32'd29862;
			35675: outdata = 32'd29861;
			35676: outdata = 32'd29860;
			35677: outdata = 32'd29859;
			35678: outdata = 32'd29858;
			35679: outdata = 32'd29857;
			35680: outdata = 32'd29856;
			35681: outdata = 32'd29855;
			35682: outdata = 32'd29854;
			35683: outdata = 32'd29853;
			35684: outdata = 32'd29852;
			35685: outdata = 32'd29851;
			35686: outdata = 32'd29850;
			35687: outdata = 32'd29849;
			35688: outdata = 32'd29848;
			35689: outdata = 32'd29847;
			35690: outdata = 32'd29846;
			35691: outdata = 32'd29845;
			35692: outdata = 32'd29844;
			35693: outdata = 32'd29843;
			35694: outdata = 32'd29842;
			35695: outdata = 32'd29841;
			35696: outdata = 32'd29840;
			35697: outdata = 32'd29839;
			35698: outdata = 32'd29838;
			35699: outdata = 32'd29837;
			35700: outdata = 32'd29836;
			35701: outdata = 32'd29835;
			35702: outdata = 32'd29834;
			35703: outdata = 32'd29833;
			35704: outdata = 32'd29832;
			35705: outdata = 32'd29831;
			35706: outdata = 32'd29830;
			35707: outdata = 32'd29829;
			35708: outdata = 32'd29828;
			35709: outdata = 32'd29827;
			35710: outdata = 32'd29826;
			35711: outdata = 32'd29825;
			35712: outdata = 32'd29824;
			35713: outdata = 32'd29823;
			35714: outdata = 32'd29822;
			35715: outdata = 32'd29821;
			35716: outdata = 32'd29820;
			35717: outdata = 32'd29819;
			35718: outdata = 32'd29818;
			35719: outdata = 32'd29817;
			35720: outdata = 32'd29816;
			35721: outdata = 32'd29815;
			35722: outdata = 32'd29814;
			35723: outdata = 32'd29813;
			35724: outdata = 32'd29812;
			35725: outdata = 32'd29811;
			35726: outdata = 32'd29810;
			35727: outdata = 32'd29809;
			35728: outdata = 32'd29808;
			35729: outdata = 32'd29807;
			35730: outdata = 32'd29806;
			35731: outdata = 32'd29805;
			35732: outdata = 32'd29804;
			35733: outdata = 32'd29803;
			35734: outdata = 32'd29802;
			35735: outdata = 32'd29801;
			35736: outdata = 32'd29800;
			35737: outdata = 32'd29799;
			35738: outdata = 32'd29798;
			35739: outdata = 32'd29797;
			35740: outdata = 32'd29796;
			35741: outdata = 32'd29795;
			35742: outdata = 32'd29794;
			35743: outdata = 32'd29793;
			35744: outdata = 32'd29792;
			35745: outdata = 32'd29791;
			35746: outdata = 32'd29790;
			35747: outdata = 32'd29789;
			35748: outdata = 32'd29788;
			35749: outdata = 32'd29787;
			35750: outdata = 32'd29786;
			35751: outdata = 32'd29785;
			35752: outdata = 32'd29784;
			35753: outdata = 32'd29783;
			35754: outdata = 32'd29782;
			35755: outdata = 32'd29781;
			35756: outdata = 32'd29780;
			35757: outdata = 32'd29779;
			35758: outdata = 32'd29778;
			35759: outdata = 32'd29777;
			35760: outdata = 32'd29776;
			35761: outdata = 32'd29775;
			35762: outdata = 32'd29774;
			35763: outdata = 32'd29773;
			35764: outdata = 32'd29772;
			35765: outdata = 32'd29771;
			35766: outdata = 32'd29770;
			35767: outdata = 32'd29769;
			35768: outdata = 32'd29768;
			35769: outdata = 32'd29767;
			35770: outdata = 32'd29766;
			35771: outdata = 32'd29765;
			35772: outdata = 32'd29764;
			35773: outdata = 32'd29763;
			35774: outdata = 32'd29762;
			35775: outdata = 32'd29761;
			35776: outdata = 32'd29760;
			35777: outdata = 32'd29759;
			35778: outdata = 32'd29758;
			35779: outdata = 32'd29757;
			35780: outdata = 32'd29756;
			35781: outdata = 32'd29755;
			35782: outdata = 32'd29754;
			35783: outdata = 32'd29753;
			35784: outdata = 32'd29752;
			35785: outdata = 32'd29751;
			35786: outdata = 32'd29750;
			35787: outdata = 32'd29749;
			35788: outdata = 32'd29748;
			35789: outdata = 32'd29747;
			35790: outdata = 32'd29746;
			35791: outdata = 32'd29745;
			35792: outdata = 32'd29744;
			35793: outdata = 32'd29743;
			35794: outdata = 32'd29742;
			35795: outdata = 32'd29741;
			35796: outdata = 32'd29740;
			35797: outdata = 32'd29739;
			35798: outdata = 32'd29738;
			35799: outdata = 32'd29737;
			35800: outdata = 32'd29736;
			35801: outdata = 32'd29735;
			35802: outdata = 32'd29734;
			35803: outdata = 32'd29733;
			35804: outdata = 32'd29732;
			35805: outdata = 32'd29731;
			35806: outdata = 32'd29730;
			35807: outdata = 32'd29729;
			35808: outdata = 32'd29728;
			35809: outdata = 32'd29727;
			35810: outdata = 32'd29726;
			35811: outdata = 32'd29725;
			35812: outdata = 32'd29724;
			35813: outdata = 32'd29723;
			35814: outdata = 32'd29722;
			35815: outdata = 32'd29721;
			35816: outdata = 32'd29720;
			35817: outdata = 32'd29719;
			35818: outdata = 32'd29718;
			35819: outdata = 32'd29717;
			35820: outdata = 32'd29716;
			35821: outdata = 32'd29715;
			35822: outdata = 32'd29714;
			35823: outdata = 32'd29713;
			35824: outdata = 32'd29712;
			35825: outdata = 32'd29711;
			35826: outdata = 32'd29710;
			35827: outdata = 32'd29709;
			35828: outdata = 32'd29708;
			35829: outdata = 32'd29707;
			35830: outdata = 32'd29706;
			35831: outdata = 32'd29705;
			35832: outdata = 32'd29704;
			35833: outdata = 32'd29703;
			35834: outdata = 32'd29702;
			35835: outdata = 32'd29701;
			35836: outdata = 32'd29700;
			35837: outdata = 32'd29699;
			35838: outdata = 32'd29698;
			35839: outdata = 32'd29697;
			35840: outdata = 32'd29696;
			35841: outdata = 32'd29695;
			35842: outdata = 32'd29694;
			35843: outdata = 32'd29693;
			35844: outdata = 32'd29692;
			35845: outdata = 32'd29691;
			35846: outdata = 32'd29690;
			35847: outdata = 32'd29689;
			35848: outdata = 32'd29688;
			35849: outdata = 32'd29687;
			35850: outdata = 32'd29686;
			35851: outdata = 32'd29685;
			35852: outdata = 32'd29684;
			35853: outdata = 32'd29683;
			35854: outdata = 32'd29682;
			35855: outdata = 32'd29681;
			35856: outdata = 32'd29680;
			35857: outdata = 32'd29679;
			35858: outdata = 32'd29678;
			35859: outdata = 32'd29677;
			35860: outdata = 32'd29676;
			35861: outdata = 32'd29675;
			35862: outdata = 32'd29674;
			35863: outdata = 32'd29673;
			35864: outdata = 32'd29672;
			35865: outdata = 32'd29671;
			35866: outdata = 32'd29670;
			35867: outdata = 32'd29669;
			35868: outdata = 32'd29668;
			35869: outdata = 32'd29667;
			35870: outdata = 32'd29666;
			35871: outdata = 32'd29665;
			35872: outdata = 32'd29664;
			35873: outdata = 32'd29663;
			35874: outdata = 32'd29662;
			35875: outdata = 32'd29661;
			35876: outdata = 32'd29660;
			35877: outdata = 32'd29659;
			35878: outdata = 32'd29658;
			35879: outdata = 32'd29657;
			35880: outdata = 32'd29656;
			35881: outdata = 32'd29655;
			35882: outdata = 32'd29654;
			35883: outdata = 32'd29653;
			35884: outdata = 32'd29652;
			35885: outdata = 32'd29651;
			35886: outdata = 32'd29650;
			35887: outdata = 32'd29649;
			35888: outdata = 32'd29648;
			35889: outdata = 32'd29647;
			35890: outdata = 32'd29646;
			35891: outdata = 32'd29645;
			35892: outdata = 32'd29644;
			35893: outdata = 32'd29643;
			35894: outdata = 32'd29642;
			35895: outdata = 32'd29641;
			35896: outdata = 32'd29640;
			35897: outdata = 32'd29639;
			35898: outdata = 32'd29638;
			35899: outdata = 32'd29637;
			35900: outdata = 32'd29636;
			35901: outdata = 32'd29635;
			35902: outdata = 32'd29634;
			35903: outdata = 32'd29633;
			35904: outdata = 32'd29632;
			35905: outdata = 32'd29631;
			35906: outdata = 32'd29630;
			35907: outdata = 32'd29629;
			35908: outdata = 32'd29628;
			35909: outdata = 32'd29627;
			35910: outdata = 32'd29626;
			35911: outdata = 32'd29625;
			35912: outdata = 32'd29624;
			35913: outdata = 32'd29623;
			35914: outdata = 32'd29622;
			35915: outdata = 32'd29621;
			35916: outdata = 32'd29620;
			35917: outdata = 32'd29619;
			35918: outdata = 32'd29618;
			35919: outdata = 32'd29617;
			35920: outdata = 32'd29616;
			35921: outdata = 32'd29615;
			35922: outdata = 32'd29614;
			35923: outdata = 32'd29613;
			35924: outdata = 32'd29612;
			35925: outdata = 32'd29611;
			35926: outdata = 32'd29610;
			35927: outdata = 32'd29609;
			35928: outdata = 32'd29608;
			35929: outdata = 32'd29607;
			35930: outdata = 32'd29606;
			35931: outdata = 32'd29605;
			35932: outdata = 32'd29604;
			35933: outdata = 32'd29603;
			35934: outdata = 32'd29602;
			35935: outdata = 32'd29601;
			35936: outdata = 32'd29600;
			35937: outdata = 32'd29599;
			35938: outdata = 32'd29598;
			35939: outdata = 32'd29597;
			35940: outdata = 32'd29596;
			35941: outdata = 32'd29595;
			35942: outdata = 32'd29594;
			35943: outdata = 32'd29593;
			35944: outdata = 32'd29592;
			35945: outdata = 32'd29591;
			35946: outdata = 32'd29590;
			35947: outdata = 32'd29589;
			35948: outdata = 32'd29588;
			35949: outdata = 32'd29587;
			35950: outdata = 32'd29586;
			35951: outdata = 32'd29585;
			35952: outdata = 32'd29584;
			35953: outdata = 32'd29583;
			35954: outdata = 32'd29582;
			35955: outdata = 32'd29581;
			35956: outdata = 32'd29580;
			35957: outdata = 32'd29579;
			35958: outdata = 32'd29578;
			35959: outdata = 32'd29577;
			35960: outdata = 32'd29576;
			35961: outdata = 32'd29575;
			35962: outdata = 32'd29574;
			35963: outdata = 32'd29573;
			35964: outdata = 32'd29572;
			35965: outdata = 32'd29571;
			35966: outdata = 32'd29570;
			35967: outdata = 32'd29569;
			35968: outdata = 32'd29568;
			35969: outdata = 32'd29567;
			35970: outdata = 32'd29566;
			35971: outdata = 32'd29565;
			35972: outdata = 32'd29564;
			35973: outdata = 32'd29563;
			35974: outdata = 32'd29562;
			35975: outdata = 32'd29561;
			35976: outdata = 32'd29560;
			35977: outdata = 32'd29559;
			35978: outdata = 32'd29558;
			35979: outdata = 32'd29557;
			35980: outdata = 32'd29556;
			35981: outdata = 32'd29555;
			35982: outdata = 32'd29554;
			35983: outdata = 32'd29553;
			35984: outdata = 32'd29552;
			35985: outdata = 32'd29551;
			35986: outdata = 32'd29550;
			35987: outdata = 32'd29549;
			35988: outdata = 32'd29548;
			35989: outdata = 32'd29547;
			35990: outdata = 32'd29546;
			35991: outdata = 32'd29545;
			35992: outdata = 32'd29544;
			35993: outdata = 32'd29543;
			35994: outdata = 32'd29542;
			35995: outdata = 32'd29541;
			35996: outdata = 32'd29540;
			35997: outdata = 32'd29539;
			35998: outdata = 32'd29538;
			35999: outdata = 32'd29537;
			36000: outdata = 32'd29536;
			36001: outdata = 32'd29535;
			36002: outdata = 32'd29534;
			36003: outdata = 32'd29533;
			36004: outdata = 32'd29532;
			36005: outdata = 32'd29531;
			36006: outdata = 32'd29530;
			36007: outdata = 32'd29529;
			36008: outdata = 32'd29528;
			36009: outdata = 32'd29527;
			36010: outdata = 32'd29526;
			36011: outdata = 32'd29525;
			36012: outdata = 32'd29524;
			36013: outdata = 32'd29523;
			36014: outdata = 32'd29522;
			36015: outdata = 32'd29521;
			36016: outdata = 32'd29520;
			36017: outdata = 32'd29519;
			36018: outdata = 32'd29518;
			36019: outdata = 32'd29517;
			36020: outdata = 32'd29516;
			36021: outdata = 32'd29515;
			36022: outdata = 32'd29514;
			36023: outdata = 32'd29513;
			36024: outdata = 32'd29512;
			36025: outdata = 32'd29511;
			36026: outdata = 32'd29510;
			36027: outdata = 32'd29509;
			36028: outdata = 32'd29508;
			36029: outdata = 32'd29507;
			36030: outdata = 32'd29506;
			36031: outdata = 32'd29505;
			36032: outdata = 32'd29504;
			36033: outdata = 32'd29503;
			36034: outdata = 32'd29502;
			36035: outdata = 32'd29501;
			36036: outdata = 32'd29500;
			36037: outdata = 32'd29499;
			36038: outdata = 32'd29498;
			36039: outdata = 32'd29497;
			36040: outdata = 32'd29496;
			36041: outdata = 32'd29495;
			36042: outdata = 32'd29494;
			36043: outdata = 32'd29493;
			36044: outdata = 32'd29492;
			36045: outdata = 32'd29491;
			36046: outdata = 32'd29490;
			36047: outdata = 32'd29489;
			36048: outdata = 32'd29488;
			36049: outdata = 32'd29487;
			36050: outdata = 32'd29486;
			36051: outdata = 32'd29485;
			36052: outdata = 32'd29484;
			36053: outdata = 32'd29483;
			36054: outdata = 32'd29482;
			36055: outdata = 32'd29481;
			36056: outdata = 32'd29480;
			36057: outdata = 32'd29479;
			36058: outdata = 32'd29478;
			36059: outdata = 32'd29477;
			36060: outdata = 32'd29476;
			36061: outdata = 32'd29475;
			36062: outdata = 32'd29474;
			36063: outdata = 32'd29473;
			36064: outdata = 32'd29472;
			36065: outdata = 32'd29471;
			36066: outdata = 32'd29470;
			36067: outdata = 32'd29469;
			36068: outdata = 32'd29468;
			36069: outdata = 32'd29467;
			36070: outdata = 32'd29466;
			36071: outdata = 32'd29465;
			36072: outdata = 32'd29464;
			36073: outdata = 32'd29463;
			36074: outdata = 32'd29462;
			36075: outdata = 32'd29461;
			36076: outdata = 32'd29460;
			36077: outdata = 32'd29459;
			36078: outdata = 32'd29458;
			36079: outdata = 32'd29457;
			36080: outdata = 32'd29456;
			36081: outdata = 32'd29455;
			36082: outdata = 32'd29454;
			36083: outdata = 32'd29453;
			36084: outdata = 32'd29452;
			36085: outdata = 32'd29451;
			36086: outdata = 32'd29450;
			36087: outdata = 32'd29449;
			36088: outdata = 32'd29448;
			36089: outdata = 32'd29447;
			36090: outdata = 32'd29446;
			36091: outdata = 32'd29445;
			36092: outdata = 32'd29444;
			36093: outdata = 32'd29443;
			36094: outdata = 32'd29442;
			36095: outdata = 32'd29441;
			36096: outdata = 32'd29440;
			36097: outdata = 32'd29439;
			36098: outdata = 32'd29438;
			36099: outdata = 32'd29437;
			36100: outdata = 32'd29436;
			36101: outdata = 32'd29435;
			36102: outdata = 32'd29434;
			36103: outdata = 32'd29433;
			36104: outdata = 32'd29432;
			36105: outdata = 32'd29431;
			36106: outdata = 32'd29430;
			36107: outdata = 32'd29429;
			36108: outdata = 32'd29428;
			36109: outdata = 32'd29427;
			36110: outdata = 32'd29426;
			36111: outdata = 32'd29425;
			36112: outdata = 32'd29424;
			36113: outdata = 32'd29423;
			36114: outdata = 32'd29422;
			36115: outdata = 32'd29421;
			36116: outdata = 32'd29420;
			36117: outdata = 32'd29419;
			36118: outdata = 32'd29418;
			36119: outdata = 32'd29417;
			36120: outdata = 32'd29416;
			36121: outdata = 32'd29415;
			36122: outdata = 32'd29414;
			36123: outdata = 32'd29413;
			36124: outdata = 32'd29412;
			36125: outdata = 32'd29411;
			36126: outdata = 32'd29410;
			36127: outdata = 32'd29409;
			36128: outdata = 32'd29408;
			36129: outdata = 32'd29407;
			36130: outdata = 32'd29406;
			36131: outdata = 32'd29405;
			36132: outdata = 32'd29404;
			36133: outdata = 32'd29403;
			36134: outdata = 32'd29402;
			36135: outdata = 32'd29401;
			36136: outdata = 32'd29400;
			36137: outdata = 32'd29399;
			36138: outdata = 32'd29398;
			36139: outdata = 32'd29397;
			36140: outdata = 32'd29396;
			36141: outdata = 32'd29395;
			36142: outdata = 32'd29394;
			36143: outdata = 32'd29393;
			36144: outdata = 32'd29392;
			36145: outdata = 32'd29391;
			36146: outdata = 32'd29390;
			36147: outdata = 32'd29389;
			36148: outdata = 32'd29388;
			36149: outdata = 32'd29387;
			36150: outdata = 32'd29386;
			36151: outdata = 32'd29385;
			36152: outdata = 32'd29384;
			36153: outdata = 32'd29383;
			36154: outdata = 32'd29382;
			36155: outdata = 32'd29381;
			36156: outdata = 32'd29380;
			36157: outdata = 32'd29379;
			36158: outdata = 32'd29378;
			36159: outdata = 32'd29377;
			36160: outdata = 32'd29376;
			36161: outdata = 32'd29375;
			36162: outdata = 32'd29374;
			36163: outdata = 32'd29373;
			36164: outdata = 32'd29372;
			36165: outdata = 32'd29371;
			36166: outdata = 32'd29370;
			36167: outdata = 32'd29369;
			36168: outdata = 32'd29368;
			36169: outdata = 32'd29367;
			36170: outdata = 32'd29366;
			36171: outdata = 32'd29365;
			36172: outdata = 32'd29364;
			36173: outdata = 32'd29363;
			36174: outdata = 32'd29362;
			36175: outdata = 32'd29361;
			36176: outdata = 32'd29360;
			36177: outdata = 32'd29359;
			36178: outdata = 32'd29358;
			36179: outdata = 32'd29357;
			36180: outdata = 32'd29356;
			36181: outdata = 32'd29355;
			36182: outdata = 32'd29354;
			36183: outdata = 32'd29353;
			36184: outdata = 32'd29352;
			36185: outdata = 32'd29351;
			36186: outdata = 32'd29350;
			36187: outdata = 32'd29349;
			36188: outdata = 32'd29348;
			36189: outdata = 32'd29347;
			36190: outdata = 32'd29346;
			36191: outdata = 32'd29345;
			36192: outdata = 32'd29344;
			36193: outdata = 32'd29343;
			36194: outdata = 32'd29342;
			36195: outdata = 32'd29341;
			36196: outdata = 32'd29340;
			36197: outdata = 32'd29339;
			36198: outdata = 32'd29338;
			36199: outdata = 32'd29337;
			36200: outdata = 32'd29336;
			36201: outdata = 32'd29335;
			36202: outdata = 32'd29334;
			36203: outdata = 32'd29333;
			36204: outdata = 32'd29332;
			36205: outdata = 32'd29331;
			36206: outdata = 32'd29330;
			36207: outdata = 32'd29329;
			36208: outdata = 32'd29328;
			36209: outdata = 32'd29327;
			36210: outdata = 32'd29326;
			36211: outdata = 32'd29325;
			36212: outdata = 32'd29324;
			36213: outdata = 32'd29323;
			36214: outdata = 32'd29322;
			36215: outdata = 32'd29321;
			36216: outdata = 32'd29320;
			36217: outdata = 32'd29319;
			36218: outdata = 32'd29318;
			36219: outdata = 32'd29317;
			36220: outdata = 32'd29316;
			36221: outdata = 32'd29315;
			36222: outdata = 32'd29314;
			36223: outdata = 32'd29313;
			36224: outdata = 32'd29312;
			36225: outdata = 32'd29311;
			36226: outdata = 32'd29310;
			36227: outdata = 32'd29309;
			36228: outdata = 32'd29308;
			36229: outdata = 32'd29307;
			36230: outdata = 32'd29306;
			36231: outdata = 32'd29305;
			36232: outdata = 32'd29304;
			36233: outdata = 32'd29303;
			36234: outdata = 32'd29302;
			36235: outdata = 32'd29301;
			36236: outdata = 32'd29300;
			36237: outdata = 32'd29299;
			36238: outdata = 32'd29298;
			36239: outdata = 32'd29297;
			36240: outdata = 32'd29296;
			36241: outdata = 32'd29295;
			36242: outdata = 32'd29294;
			36243: outdata = 32'd29293;
			36244: outdata = 32'd29292;
			36245: outdata = 32'd29291;
			36246: outdata = 32'd29290;
			36247: outdata = 32'd29289;
			36248: outdata = 32'd29288;
			36249: outdata = 32'd29287;
			36250: outdata = 32'd29286;
			36251: outdata = 32'd29285;
			36252: outdata = 32'd29284;
			36253: outdata = 32'd29283;
			36254: outdata = 32'd29282;
			36255: outdata = 32'd29281;
			36256: outdata = 32'd29280;
			36257: outdata = 32'd29279;
			36258: outdata = 32'd29278;
			36259: outdata = 32'd29277;
			36260: outdata = 32'd29276;
			36261: outdata = 32'd29275;
			36262: outdata = 32'd29274;
			36263: outdata = 32'd29273;
			36264: outdata = 32'd29272;
			36265: outdata = 32'd29271;
			36266: outdata = 32'd29270;
			36267: outdata = 32'd29269;
			36268: outdata = 32'd29268;
			36269: outdata = 32'd29267;
			36270: outdata = 32'd29266;
			36271: outdata = 32'd29265;
			36272: outdata = 32'd29264;
			36273: outdata = 32'd29263;
			36274: outdata = 32'd29262;
			36275: outdata = 32'd29261;
			36276: outdata = 32'd29260;
			36277: outdata = 32'd29259;
			36278: outdata = 32'd29258;
			36279: outdata = 32'd29257;
			36280: outdata = 32'd29256;
			36281: outdata = 32'd29255;
			36282: outdata = 32'd29254;
			36283: outdata = 32'd29253;
			36284: outdata = 32'd29252;
			36285: outdata = 32'd29251;
			36286: outdata = 32'd29250;
			36287: outdata = 32'd29249;
			36288: outdata = 32'd29248;
			36289: outdata = 32'd29247;
			36290: outdata = 32'd29246;
			36291: outdata = 32'd29245;
			36292: outdata = 32'd29244;
			36293: outdata = 32'd29243;
			36294: outdata = 32'd29242;
			36295: outdata = 32'd29241;
			36296: outdata = 32'd29240;
			36297: outdata = 32'd29239;
			36298: outdata = 32'd29238;
			36299: outdata = 32'd29237;
			36300: outdata = 32'd29236;
			36301: outdata = 32'd29235;
			36302: outdata = 32'd29234;
			36303: outdata = 32'd29233;
			36304: outdata = 32'd29232;
			36305: outdata = 32'd29231;
			36306: outdata = 32'd29230;
			36307: outdata = 32'd29229;
			36308: outdata = 32'd29228;
			36309: outdata = 32'd29227;
			36310: outdata = 32'd29226;
			36311: outdata = 32'd29225;
			36312: outdata = 32'd29224;
			36313: outdata = 32'd29223;
			36314: outdata = 32'd29222;
			36315: outdata = 32'd29221;
			36316: outdata = 32'd29220;
			36317: outdata = 32'd29219;
			36318: outdata = 32'd29218;
			36319: outdata = 32'd29217;
			36320: outdata = 32'd29216;
			36321: outdata = 32'd29215;
			36322: outdata = 32'd29214;
			36323: outdata = 32'd29213;
			36324: outdata = 32'd29212;
			36325: outdata = 32'd29211;
			36326: outdata = 32'd29210;
			36327: outdata = 32'd29209;
			36328: outdata = 32'd29208;
			36329: outdata = 32'd29207;
			36330: outdata = 32'd29206;
			36331: outdata = 32'd29205;
			36332: outdata = 32'd29204;
			36333: outdata = 32'd29203;
			36334: outdata = 32'd29202;
			36335: outdata = 32'd29201;
			36336: outdata = 32'd29200;
			36337: outdata = 32'd29199;
			36338: outdata = 32'd29198;
			36339: outdata = 32'd29197;
			36340: outdata = 32'd29196;
			36341: outdata = 32'd29195;
			36342: outdata = 32'd29194;
			36343: outdata = 32'd29193;
			36344: outdata = 32'd29192;
			36345: outdata = 32'd29191;
			36346: outdata = 32'd29190;
			36347: outdata = 32'd29189;
			36348: outdata = 32'd29188;
			36349: outdata = 32'd29187;
			36350: outdata = 32'd29186;
			36351: outdata = 32'd29185;
			36352: outdata = 32'd29184;
			36353: outdata = 32'd29183;
			36354: outdata = 32'd29182;
			36355: outdata = 32'd29181;
			36356: outdata = 32'd29180;
			36357: outdata = 32'd29179;
			36358: outdata = 32'd29178;
			36359: outdata = 32'd29177;
			36360: outdata = 32'd29176;
			36361: outdata = 32'd29175;
			36362: outdata = 32'd29174;
			36363: outdata = 32'd29173;
			36364: outdata = 32'd29172;
			36365: outdata = 32'd29171;
			36366: outdata = 32'd29170;
			36367: outdata = 32'd29169;
			36368: outdata = 32'd29168;
			36369: outdata = 32'd29167;
			36370: outdata = 32'd29166;
			36371: outdata = 32'd29165;
			36372: outdata = 32'd29164;
			36373: outdata = 32'd29163;
			36374: outdata = 32'd29162;
			36375: outdata = 32'd29161;
			36376: outdata = 32'd29160;
			36377: outdata = 32'd29159;
			36378: outdata = 32'd29158;
			36379: outdata = 32'd29157;
			36380: outdata = 32'd29156;
			36381: outdata = 32'd29155;
			36382: outdata = 32'd29154;
			36383: outdata = 32'd29153;
			36384: outdata = 32'd29152;
			36385: outdata = 32'd29151;
			36386: outdata = 32'd29150;
			36387: outdata = 32'd29149;
			36388: outdata = 32'd29148;
			36389: outdata = 32'd29147;
			36390: outdata = 32'd29146;
			36391: outdata = 32'd29145;
			36392: outdata = 32'd29144;
			36393: outdata = 32'd29143;
			36394: outdata = 32'd29142;
			36395: outdata = 32'd29141;
			36396: outdata = 32'd29140;
			36397: outdata = 32'd29139;
			36398: outdata = 32'd29138;
			36399: outdata = 32'd29137;
			36400: outdata = 32'd29136;
			36401: outdata = 32'd29135;
			36402: outdata = 32'd29134;
			36403: outdata = 32'd29133;
			36404: outdata = 32'd29132;
			36405: outdata = 32'd29131;
			36406: outdata = 32'd29130;
			36407: outdata = 32'd29129;
			36408: outdata = 32'd29128;
			36409: outdata = 32'd29127;
			36410: outdata = 32'd29126;
			36411: outdata = 32'd29125;
			36412: outdata = 32'd29124;
			36413: outdata = 32'd29123;
			36414: outdata = 32'd29122;
			36415: outdata = 32'd29121;
			36416: outdata = 32'd29120;
			36417: outdata = 32'd29119;
			36418: outdata = 32'd29118;
			36419: outdata = 32'd29117;
			36420: outdata = 32'd29116;
			36421: outdata = 32'd29115;
			36422: outdata = 32'd29114;
			36423: outdata = 32'd29113;
			36424: outdata = 32'd29112;
			36425: outdata = 32'd29111;
			36426: outdata = 32'd29110;
			36427: outdata = 32'd29109;
			36428: outdata = 32'd29108;
			36429: outdata = 32'd29107;
			36430: outdata = 32'd29106;
			36431: outdata = 32'd29105;
			36432: outdata = 32'd29104;
			36433: outdata = 32'd29103;
			36434: outdata = 32'd29102;
			36435: outdata = 32'd29101;
			36436: outdata = 32'd29100;
			36437: outdata = 32'd29099;
			36438: outdata = 32'd29098;
			36439: outdata = 32'd29097;
			36440: outdata = 32'd29096;
			36441: outdata = 32'd29095;
			36442: outdata = 32'd29094;
			36443: outdata = 32'd29093;
			36444: outdata = 32'd29092;
			36445: outdata = 32'd29091;
			36446: outdata = 32'd29090;
			36447: outdata = 32'd29089;
			36448: outdata = 32'd29088;
			36449: outdata = 32'd29087;
			36450: outdata = 32'd29086;
			36451: outdata = 32'd29085;
			36452: outdata = 32'd29084;
			36453: outdata = 32'd29083;
			36454: outdata = 32'd29082;
			36455: outdata = 32'd29081;
			36456: outdata = 32'd29080;
			36457: outdata = 32'd29079;
			36458: outdata = 32'd29078;
			36459: outdata = 32'd29077;
			36460: outdata = 32'd29076;
			36461: outdata = 32'd29075;
			36462: outdata = 32'd29074;
			36463: outdata = 32'd29073;
			36464: outdata = 32'd29072;
			36465: outdata = 32'd29071;
			36466: outdata = 32'd29070;
			36467: outdata = 32'd29069;
			36468: outdata = 32'd29068;
			36469: outdata = 32'd29067;
			36470: outdata = 32'd29066;
			36471: outdata = 32'd29065;
			36472: outdata = 32'd29064;
			36473: outdata = 32'd29063;
			36474: outdata = 32'd29062;
			36475: outdata = 32'd29061;
			36476: outdata = 32'd29060;
			36477: outdata = 32'd29059;
			36478: outdata = 32'd29058;
			36479: outdata = 32'd29057;
			36480: outdata = 32'd29056;
			36481: outdata = 32'd29055;
			36482: outdata = 32'd29054;
			36483: outdata = 32'd29053;
			36484: outdata = 32'd29052;
			36485: outdata = 32'd29051;
			36486: outdata = 32'd29050;
			36487: outdata = 32'd29049;
			36488: outdata = 32'd29048;
			36489: outdata = 32'd29047;
			36490: outdata = 32'd29046;
			36491: outdata = 32'd29045;
			36492: outdata = 32'd29044;
			36493: outdata = 32'd29043;
			36494: outdata = 32'd29042;
			36495: outdata = 32'd29041;
			36496: outdata = 32'd29040;
			36497: outdata = 32'd29039;
			36498: outdata = 32'd29038;
			36499: outdata = 32'd29037;
			36500: outdata = 32'd29036;
			36501: outdata = 32'd29035;
			36502: outdata = 32'd29034;
			36503: outdata = 32'd29033;
			36504: outdata = 32'd29032;
			36505: outdata = 32'd29031;
			36506: outdata = 32'd29030;
			36507: outdata = 32'd29029;
			36508: outdata = 32'd29028;
			36509: outdata = 32'd29027;
			36510: outdata = 32'd29026;
			36511: outdata = 32'd29025;
			36512: outdata = 32'd29024;
			36513: outdata = 32'd29023;
			36514: outdata = 32'd29022;
			36515: outdata = 32'd29021;
			36516: outdata = 32'd29020;
			36517: outdata = 32'd29019;
			36518: outdata = 32'd29018;
			36519: outdata = 32'd29017;
			36520: outdata = 32'd29016;
			36521: outdata = 32'd29015;
			36522: outdata = 32'd29014;
			36523: outdata = 32'd29013;
			36524: outdata = 32'd29012;
			36525: outdata = 32'd29011;
			36526: outdata = 32'd29010;
			36527: outdata = 32'd29009;
			36528: outdata = 32'd29008;
			36529: outdata = 32'd29007;
			36530: outdata = 32'd29006;
			36531: outdata = 32'd29005;
			36532: outdata = 32'd29004;
			36533: outdata = 32'd29003;
			36534: outdata = 32'd29002;
			36535: outdata = 32'd29001;
			36536: outdata = 32'd29000;
			36537: outdata = 32'd28999;
			36538: outdata = 32'd28998;
			36539: outdata = 32'd28997;
			36540: outdata = 32'd28996;
			36541: outdata = 32'd28995;
			36542: outdata = 32'd28994;
			36543: outdata = 32'd28993;
			36544: outdata = 32'd28992;
			36545: outdata = 32'd28991;
			36546: outdata = 32'd28990;
			36547: outdata = 32'd28989;
			36548: outdata = 32'd28988;
			36549: outdata = 32'd28987;
			36550: outdata = 32'd28986;
			36551: outdata = 32'd28985;
			36552: outdata = 32'd28984;
			36553: outdata = 32'd28983;
			36554: outdata = 32'd28982;
			36555: outdata = 32'd28981;
			36556: outdata = 32'd28980;
			36557: outdata = 32'd28979;
			36558: outdata = 32'd28978;
			36559: outdata = 32'd28977;
			36560: outdata = 32'd28976;
			36561: outdata = 32'd28975;
			36562: outdata = 32'd28974;
			36563: outdata = 32'd28973;
			36564: outdata = 32'd28972;
			36565: outdata = 32'd28971;
			36566: outdata = 32'd28970;
			36567: outdata = 32'd28969;
			36568: outdata = 32'd28968;
			36569: outdata = 32'd28967;
			36570: outdata = 32'd28966;
			36571: outdata = 32'd28965;
			36572: outdata = 32'd28964;
			36573: outdata = 32'd28963;
			36574: outdata = 32'd28962;
			36575: outdata = 32'd28961;
			36576: outdata = 32'd28960;
			36577: outdata = 32'd28959;
			36578: outdata = 32'd28958;
			36579: outdata = 32'd28957;
			36580: outdata = 32'd28956;
			36581: outdata = 32'd28955;
			36582: outdata = 32'd28954;
			36583: outdata = 32'd28953;
			36584: outdata = 32'd28952;
			36585: outdata = 32'd28951;
			36586: outdata = 32'd28950;
			36587: outdata = 32'd28949;
			36588: outdata = 32'd28948;
			36589: outdata = 32'd28947;
			36590: outdata = 32'd28946;
			36591: outdata = 32'd28945;
			36592: outdata = 32'd28944;
			36593: outdata = 32'd28943;
			36594: outdata = 32'd28942;
			36595: outdata = 32'd28941;
			36596: outdata = 32'd28940;
			36597: outdata = 32'd28939;
			36598: outdata = 32'd28938;
			36599: outdata = 32'd28937;
			36600: outdata = 32'd28936;
			36601: outdata = 32'd28935;
			36602: outdata = 32'd28934;
			36603: outdata = 32'd28933;
			36604: outdata = 32'd28932;
			36605: outdata = 32'd28931;
			36606: outdata = 32'd28930;
			36607: outdata = 32'd28929;
			36608: outdata = 32'd28928;
			36609: outdata = 32'd28927;
			36610: outdata = 32'd28926;
			36611: outdata = 32'd28925;
			36612: outdata = 32'd28924;
			36613: outdata = 32'd28923;
			36614: outdata = 32'd28922;
			36615: outdata = 32'd28921;
			36616: outdata = 32'd28920;
			36617: outdata = 32'd28919;
			36618: outdata = 32'd28918;
			36619: outdata = 32'd28917;
			36620: outdata = 32'd28916;
			36621: outdata = 32'd28915;
			36622: outdata = 32'd28914;
			36623: outdata = 32'd28913;
			36624: outdata = 32'd28912;
			36625: outdata = 32'd28911;
			36626: outdata = 32'd28910;
			36627: outdata = 32'd28909;
			36628: outdata = 32'd28908;
			36629: outdata = 32'd28907;
			36630: outdata = 32'd28906;
			36631: outdata = 32'd28905;
			36632: outdata = 32'd28904;
			36633: outdata = 32'd28903;
			36634: outdata = 32'd28902;
			36635: outdata = 32'd28901;
			36636: outdata = 32'd28900;
			36637: outdata = 32'd28899;
			36638: outdata = 32'd28898;
			36639: outdata = 32'd28897;
			36640: outdata = 32'd28896;
			36641: outdata = 32'd28895;
			36642: outdata = 32'd28894;
			36643: outdata = 32'd28893;
			36644: outdata = 32'd28892;
			36645: outdata = 32'd28891;
			36646: outdata = 32'd28890;
			36647: outdata = 32'd28889;
			36648: outdata = 32'd28888;
			36649: outdata = 32'd28887;
			36650: outdata = 32'd28886;
			36651: outdata = 32'd28885;
			36652: outdata = 32'd28884;
			36653: outdata = 32'd28883;
			36654: outdata = 32'd28882;
			36655: outdata = 32'd28881;
			36656: outdata = 32'd28880;
			36657: outdata = 32'd28879;
			36658: outdata = 32'd28878;
			36659: outdata = 32'd28877;
			36660: outdata = 32'd28876;
			36661: outdata = 32'd28875;
			36662: outdata = 32'd28874;
			36663: outdata = 32'd28873;
			36664: outdata = 32'd28872;
			36665: outdata = 32'd28871;
			36666: outdata = 32'd28870;
			36667: outdata = 32'd28869;
			36668: outdata = 32'd28868;
			36669: outdata = 32'd28867;
			36670: outdata = 32'd28866;
			36671: outdata = 32'd28865;
			36672: outdata = 32'd28864;
			36673: outdata = 32'd28863;
			36674: outdata = 32'd28862;
			36675: outdata = 32'd28861;
			36676: outdata = 32'd28860;
			36677: outdata = 32'd28859;
			36678: outdata = 32'd28858;
			36679: outdata = 32'd28857;
			36680: outdata = 32'd28856;
			36681: outdata = 32'd28855;
			36682: outdata = 32'd28854;
			36683: outdata = 32'd28853;
			36684: outdata = 32'd28852;
			36685: outdata = 32'd28851;
			36686: outdata = 32'd28850;
			36687: outdata = 32'd28849;
			36688: outdata = 32'd28848;
			36689: outdata = 32'd28847;
			36690: outdata = 32'd28846;
			36691: outdata = 32'd28845;
			36692: outdata = 32'd28844;
			36693: outdata = 32'd28843;
			36694: outdata = 32'd28842;
			36695: outdata = 32'd28841;
			36696: outdata = 32'd28840;
			36697: outdata = 32'd28839;
			36698: outdata = 32'd28838;
			36699: outdata = 32'd28837;
			36700: outdata = 32'd28836;
			36701: outdata = 32'd28835;
			36702: outdata = 32'd28834;
			36703: outdata = 32'd28833;
			36704: outdata = 32'd28832;
			36705: outdata = 32'd28831;
			36706: outdata = 32'd28830;
			36707: outdata = 32'd28829;
			36708: outdata = 32'd28828;
			36709: outdata = 32'd28827;
			36710: outdata = 32'd28826;
			36711: outdata = 32'd28825;
			36712: outdata = 32'd28824;
			36713: outdata = 32'd28823;
			36714: outdata = 32'd28822;
			36715: outdata = 32'd28821;
			36716: outdata = 32'd28820;
			36717: outdata = 32'd28819;
			36718: outdata = 32'd28818;
			36719: outdata = 32'd28817;
			36720: outdata = 32'd28816;
			36721: outdata = 32'd28815;
			36722: outdata = 32'd28814;
			36723: outdata = 32'd28813;
			36724: outdata = 32'd28812;
			36725: outdata = 32'd28811;
			36726: outdata = 32'd28810;
			36727: outdata = 32'd28809;
			36728: outdata = 32'd28808;
			36729: outdata = 32'd28807;
			36730: outdata = 32'd28806;
			36731: outdata = 32'd28805;
			36732: outdata = 32'd28804;
			36733: outdata = 32'd28803;
			36734: outdata = 32'd28802;
			36735: outdata = 32'd28801;
			36736: outdata = 32'd28800;
			36737: outdata = 32'd28799;
			36738: outdata = 32'd28798;
			36739: outdata = 32'd28797;
			36740: outdata = 32'd28796;
			36741: outdata = 32'd28795;
			36742: outdata = 32'd28794;
			36743: outdata = 32'd28793;
			36744: outdata = 32'd28792;
			36745: outdata = 32'd28791;
			36746: outdata = 32'd28790;
			36747: outdata = 32'd28789;
			36748: outdata = 32'd28788;
			36749: outdata = 32'd28787;
			36750: outdata = 32'd28786;
			36751: outdata = 32'd28785;
			36752: outdata = 32'd28784;
			36753: outdata = 32'd28783;
			36754: outdata = 32'd28782;
			36755: outdata = 32'd28781;
			36756: outdata = 32'd28780;
			36757: outdata = 32'd28779;
			36758: outdata = 32'd28778;
			36759: outdata = 32'd28777;
			36760: outdata = 32'd28776;
			36761: outdata = 32'd28775;
			36762: outdata = 32'd28774;
			36763: outdata = 32'd28773;
			36764: outdata = 32'd28772;
			36765: outdata = 32'd28771;
			36766: outdata = 32'd28770;
			36767: outdata = 32'd28769;
			36768: outdata = 32'd28768;
			36769: outdata = 32'd28767;
			36770: outdata = 32'd28766;
			36771: outdata = 32'd28765;
			36772: outdata = 32'd28764;
			36773: outdata = 32'd28763;
			36774: outdata = 32'd28762;
			36775: outdata = 32'd28761;
			36776: outdata = 32'd28760;
			36777: outdata = 32'd28759;
			36778: outdata = 32'd28758;
			36779: outdata = 32'd28757;
			36780: outdata = 32'd28756;
			36781: outdata = 32'd28755;
			36782: outdata = 32'd28754;
			36783: outdata = 32'd28753;
			36784: outdata = 32'd28752;
			36785: outdata = 32'd28751;
			36786: outdata = 32'd28750;
			36787: outdata = 32'd28749;
			36788: outdata = 32'd28748;
			36789: outdata = 32'd28747;
			36790: outdata = 32'd28746;
			36791: outdata = 32'd28745;
			36792: outdata = 32'd28744;
			36793: outdata = 32'd28743;
			36794: outdata = 32'd28742;
			36795: outdata = 32'd28741;
			36796: outdata = 32'd28740;
			36797: outdata = 32'd28739;
			36798: outdata = 32'd28738;
			36799: outdata = 32'd28737;
			36800: outdata = 32'd28736;
			36801: outdata = 32'd28735;
			36802: outdata = 32'd28734;
			36803: outdata = 32'd28733;
			36804: outdata = 32'd28732;
			36805: outdata = 32'd28731;
			36806: outdata = 32'd28730;
			36807: outdata = 32'd28729;
			36808: outdata = 32'd28728;
			36809: outdata = 32'd28727;
			36810: outdata = 32'd28726;
			36811: outdata = 32'd28725;
			36812: outdata = 32'd28724;
			36813: outdata = 32'd28723;
			36814: outdata = 32'd28722;
			36815: outdata = 32'd28721;
			36816: outdata = 32'd28720;
			36817: outdata = 32'd28719;
			36818: outdata = 32'd28718;
			36819: outdata = 32'd28717;
			36820: outdata = 32'd28716;
			36821: outdata = 32'd28715;
			36822: outdata = 32'd28714;
			36823: outdata = 32'd28713;
			36824: outdata = 32'd28712;
			36825: outdata = 32'd28711;
			36826: outdata = 32'd28710;
			36827: outdata = 32'd28709;
			36828: outdata = 32'd28708;
			36829: outdata = 32'd28707;
			36830: outdata = 32'd28706;
			36831: outdata = 32'd28705;
			36832: outdata = 32'd28704;
			36833: outdata = 32'd28703;
			36834: outdata = 32'd28702;
			36835: outdata = 32'd28701;
			36836: outdata = 32'd28700;
			36837: outdata = 32'd28699;
			36838: outdata = 32'd28698;
			36839: outdata = 32'd28697;
			36840: outdata = 32'd28696;
			36841: outdata = 32'd28695;
			36842: outdata = 32'd28694;
			36843: outdata = 32'd28693;
			36844: outdata = 32'd28692;
			36845: outdata = 32'd28691;
			36846: outdata = 32'd28690;
			36847: outdata = 32'd28689;
			36848: outdata = 32'd28688;
			36849: outdata = 32'd28687;
			36850: outdata = 32'd28686;
			36851: outdata = 32'd28685;
			36852: outdata = 32'd28684;
			36853: outdata = 32'd28683;
			36854: outdata = 32'd28682;
			36855: outdata = 32'd28681;
			36856: outdata = 32'd28680;
			36857: outdata = 32'd28679;
			36858: outdata = 32'd28678;
			36859: outdata = 32'd28677;
			36860: outdata = 32'd28676;
			36861: outdata = 32'd28675;
			36862: outdata = 32'd28674;
			36863: outdata = 32'd28673;
			36864: outdata = 32'd28672;
			36865: outdata = 32'd28671;
			36866: outdata = 32'd28670;
			36867: outdata = 32'd28669;
			36868: outdata = 32'd28668;
			36869: outdata = 32'd28667;
			36870: outdata = 32'd28666;
			36871: outdata = 32'd28665;
			36872: outdata = 32'd28664;
			36873: outdata = 32'd28663;
			36874: outdata = 32'd28662;
			36875: outdata = 32'd28661;
			36876: outdata = 32'd28660;
			36877: outdata = 32'd28659;
			36878: outdata = 32'd28658;
			36879: outdata = 32'd28657;
			36880: outdata = 32'd28656;
			36881: outdata = 32'd28655;
			36882: outdata = 32'd28654;
			36883: outdata = 32'd28653;
			36884: outdata = 32'd28652;
			36885: outdata = 32'd28651;
			36886: outdata = 32'd28650;
			36887: outdata = 32'd28649;
			36888: outdata = 32'd28648;
			36889: outdata = 32'd28647;
			36890: outdata = 32'd28646;
			36891: outdata = 32'd28645;
			36892: outdata = 32'd28644;
			36893: outdata = 32'd28643;
			36894: outdata = 32'd28642;
			36895: outdata = 32'd28641;
			36896: outdata = 32'd28640;
			36897: outdata = 32'd28639;
			36898: outdata = 32'd28638;
			36899: outdata = 32'd28637;
			36900: outdata = 32'd28636;
			36901: outdata = 32'd28635;
			36902: outdata = 32'd28634;
			36903: outdata = 32'd28633;
			36904: outdata = 32'd28632;
			36905: outdata = 32'd28631;
			36906: outdata = 32'd28630;
			36907: outdata = 32'd28629;
			36908: outdata = 32'd28628;
			36909: outdata = 32'd28627;
			36910: outdata = 32'd28626;
			36911: outdata = 32'd28625;
			36912: outdata = 32'd28624;
			36913: outdata = 32'd28623;
			36914: outdata = 32'd28622;
			36915: outdata = 32'd28621;
			36916: outdata = 32'd28620;
			36917: outdata = 32'd28619;
			36918: outdata = 32'd28618;
			36919: outdata = 32'd28617;
			36920: outdata = 32'd28616;
			36921: outdata = 32'd28615;
			36922: outdata = 32'd28614;
			36923: outdata = 32'd28613;
			36924: outdata = 32'd28612;
			36925: outdata = 32'd28611;
			36926: outdata = 32'd28610;
			36927: outdata = 32'd28609;
			36928: outdata = 32'd28608;
			36929: outdata = 32'd28607;
			36930: outdata = 32'd28606;
			36931: outdata = 32'd28605;
			36932: outdata = 32'd28604;
			36933: outdata = 32'd28603;
			36934: outdata = 32'd28602;
			36935: outdata = 32'd28601;
			36936: outdata = 32'd28600;
			36937: outdata = 32'd28599;
			36938: outdata = 32'd28598;
			36939: outdata = 32'd28597;
			36940: outdata = 32'd28596;
			36941: outdata = 32'd28595;
			36942: outdata = 32'd28594;
			36943: outdata = 32'd28593;
			36944: outdata = 32'd28592;
			36945: outdata = 32'd28591;
			36946: outdata = 32'd28590;
			36947: outdata = 32'd28589;
			36948: outdata = 32'd28588;
			36949: outdata = 32'd28587;
			36950: outdata = 32'd28586;
			36951: outdata = 32'd28585;
			36952: outdata = 32'd28584;
			36953: outdata = 32'd28583;
			36954: outdata = 32'd28582;
			36955: outdata = 32'd28581;
			36956: outdata = 32'd28580;
			36957: outdata = 32'd28579;
			36958: outdata = 32'd28578;
			36959: outdata = 32'd28577;
			36960: outdata = 32'd28576;
			36961: outdata = 32'd28575;
			36962: outdata = 32'd28574;
			36963: outdata = 32'd28573;
			36964: outdata = 32'd28572;
			36965: outdata = 32'd28571;
			36966: outdata = 32'd28570;
			36967: outdata = 32'd28569;
			36968: outdata = 32'd28568;
			36969: outdata = 32'd28567;
			36970: outdata = 32'd28566;
			36971: outdata = 32'd28565;
			36972: outdata = 32'd28564;
			36973: outdata = 32'd28563;
			36974: outdata = 32'd28562;
			36975: outdata = 32'd28561;
			36976: outdata = 32'd28560;
			36977: outdata = 32'd28559;
			36978: outdata = 32'd28558;
			36979: outdata = 32'd28557;
			36980: outdata = 32'd28556;
			36981: outdata = 32'd28555;
			36982: outdata = 32'd28554;
			36983: outdata = 32'd28553;
			36984: outdata = 32'd28552;
			36985: outdata = 32'd28551;
			36986: outdata = 32'd28550;
			36987: outdata = 32'd28549;
			36988: outdata = 32'd28548;
			36989: outdata = 32'd28547;
			36990: outdata = 32'd28546;
			36991: outdata = 32'd28545;
			36992: outdata = 32'd28544;
			36993: outdata = 32'd28543;
			36994: outdata = 32'd28542;
			36995: outdata = 32'd28541;
			36996: outdata = 32'd28540;
			36997: outdata = 32'd28539;
			36998: outdata = 32'd28538;
			36999: outdata = 32'd28537;
			37000: outdata = 32'd28536;
			37001: outdata = 32'd28535;
			37002: outdata = 32'd28534;
			37003: outdata = 32'd28533;
			37004: outdata = 32'd28532;
			37005: outdata = 32'd28531;
			37006: outdata = 32'd28530;
			37007: outdata = 32'd28529;
			37008: outdata = 32'd28528;
			37009: outdata = 32'd28527;
			37010: outdata = 32'd28526;
			37011: outdata = 32'd28525;
			37012: outdata = 32'd28524;
			37013: outdata = 32'd28523;
			37014: outdata = 32'd28522;
			37015: outdata = 32'd28521;
			37016: outdata = 32'd28520;
			37017: outdata = 32'd28519;
			37018: outdata = 32'd28518;
			37019: outdata = 32'd28517;
			37020: outdata = 32'd28516;
			37021: outdata = 32'd28515;
			37022: outdata = 32'd28514;
			37023: outdata = 32'd28513;
			37024: outdata = 32'd28512;
			37025: outdata = 32'd28511;
			37026: outdata = 32'd28510;
			37027: outdata = 32'd28509;
			37028: outdata = 32'd28508;
			37029: outdata = 32'd28507;
			37030: outdata = 32'd28506;
			37031: outdata = 32'd28505;
			37032: outdata = 32'd28504;
			37033: outdata = 32'd28503;
			37034: outdata = 32'd28502;
			37035: outdata = 32'd28501;
			37036: outdata = 32'd28500;
			37037: outdata = 32'd28499;
			37038: outdata = 32'd28498;
			37039: outdata = 32'd28497;
			37040: outdata = 32'd28496;
			37041: outdata = 32'd28495;
			37042: outdata = 32'd28494;
			37043: outdata = 32'd28493;
			37044: outdata = 32'd28492;
			37045: outdata = 32'd28491;
			37046: outdata = 32'd28490;
			37047: outdata = 32'd28489;
			37048: outdata = 32'd28488;
			37049: outdata = 32'd28487;
			37050: outdata = 32'd28486;
			37051: outdata = 32'd28485;
			37052: outdata = 32'd28484;
			37053: outdata = 32'd28483;
			37054: outdata = 32'd28482;
			37055: outdata = 32'd28481;
			37056: outdata = 32'd28480;
			37057: outdata = 32'd28479;
			37058: outdata = 32'd28478;
			37059: outdata = 32'd28477;
			37060: outdata = 32'd28476;
			37061: outdata = 32'd28475;
			37062: outdata = 32'd28474;
			37063: outdata = 32'd28473;
			37064: outdata = 32'd28472;
			37065: outdata = 32'd28471;
			37066: outdata = 32'd28470;
			37067: outdata = 32'd28469;
			37068: outdata = 32'd28468;
			37069: outdata = 32'd28467;
			37070: outdata = 32'd28466;
			37071: outdata = 32'd28465;
			37072: outdata = 32'd28464;
			37073: outdata = 32'd28463;
			37074: outdata = 32'd28462;
			37075: outdata = 32'd28461;
			37076: outdata = 32'd28460;
			37077: outdata = 32'd28459;
			37078: outdata = 32'd28458;
			37079: outdata = 32'd28457;
			37080: outdata = 32'd28456;
			37081: outdata = 32'd28455;
			37082: outdata = 32'd28454;
			37083: outdata = 32'd28453;
			37084: outdata = 32'd28452;
			37085: outdata = 32'd28451;
			37086: outdata = 32'd28450;
			37087: outdata = 32'd28449;
			37088: outdata = 32'd28448;
			37089: outdata = 32'd28447;
			37090: outdata = 32'd28446;
			37091: outdata = 32'd28445;
			37092: outdata = 32'd28444;
			37093: outdata = 32'd28443;
			37094: outdata = 32'd28442;
			37095: outdata = 32'd28441;
			37096: outdata = 32'd28440;
			37097: outdata = 32'd28439;
			37098: outdata = 32'd28438;
			37099: outdata = 32'd28437;
			37100: outdata = 32'd28436;
			37101: outdata = 32'd28435;
			37102: outdata = 32'd28434;
			37103: outdata = 32'd28433;
			37104: outdata = 32'd28432;
			37105: outdata = 32'd28431;
			37106: outdata = 32'd28430;
			37107: outdata = 32'd28429;
			37108: outdata = 32'd28428;
			37109: outdata = 32'd28427;
			37110: outdata = 32'd28426;
			37111: outdata = 32'd28425;
			37112: outdata = 32'd28424;
			37113: outdata = 32'd28423;
			37114: outdata = 32'd28422;
			37115: outdata = 32'd28421;
			37116: outdata = 32'd28420;
			37117: outdata = 32'd28419;
			37118: outdata = 32'd28418;
			37119: outdata = 32'd28417;
			37120: outdata = 32'd28416;
			37121: outdata = 32'd28415;
			37122: outdata = 32'd28414;
			37123: outdata = 32'd28413;
			37124: outdata = 32'd28412;
			37125: outdata = 32'd28411;
			37126: outdata = 32'd28410;
			37127: outdata = 32'd28409;
			37128: outdata = 32'd28408;
			37129: outdata = 32'd28407;
			37130: outdata = 32'd28406;
			37131: outdata = 32'd28405;
			37132: outdata = 32'd28404;
			37133: outdata = 32'd28403;
			37134: outdata = 32'd28402;
			37135: outdata = 32'd28401;
			37136: outdata = 32'd28400;
			37137: outdata = 32'd28399;
			37138: outdata = 32'd28398;
			37139: outdata = 32'd28397;
			37140: outdata = 32'd28396;
			37141: outdata = 32'd28395;
			37142: outdata = 32'd28394;
			37143: outdata = 32'd28393;
			37144: outdata = 32'd28392;
			37145: outdata = 32'd28391;
			37146: outdata = 32'd28390;
			37147: outdata = 32'd28389;
			37148: outdata = 32'd28388;
			37149: outdata = 32'd28387;
			37150: outdata = 32'd28386;
			37151: outdata = 32'd28385;
			37152: outdata = 32'd28384;
			37153: outdata = 32'd28383;
			37154: outdata = 32'd28382;
			37155: outdata = 32'd28381;
			37156: outdata = 32'd28380;
			37157: outdata = 32'd28379;
			37158: outdata = 32'd28378;
			37159: outdata = 32'd28377;
			37160: outdata = 32'd28376;
			37161: outdata = 32'd28375;
			37162: outdata = 32'd28374;
			37163: outdata = 32'd28373;
			37164: outdata = 32'd28372;
			37165: outdata = 32'd28371;
			37166: outdata = 32'd28370;
			37167: outdata = 32'd28369;
			37168: outdata = 32'd28368;
			37169: outdata = 32'd28367;
			37170: outdata = 32'd28366;
			37171: outdata = 32'd28365;
			37172: outdata = 32'd28364;
			37173: outdata = 32'd28363;
			37174: outdata = 32'd28362;
			37175: outdata = 32'd28361;
			37176: outdata = 32'd28360;
			37177: outdata = 32'd28359;
			37178: outdata = 32'd28358;
			37179: outdata = 32'd28357;
			37180: outdata = 32'd28356;
			37181: outdata = 32'd28355;
			37182: outdata = 32'd28354;
			37183: outdata = 32'd28353;
			37184: outdata = 32'd28352;
			37185: outdata = 32'd28351;
			37186: outdata = 32'd28350;
			37187: outdata = 32'd28349;
			37188: outdata = 32'd28348;
			37189: outdata = 32'd28347;
			37190: outdata = 32'd28346;
			37191: outdata = 32'd28345;
			37192: outdata = 32'd28344;
			37193: outdata = 32'd28343;
			37194: outdata = 32'd28342;
			37195: outdata = 32'd28341;
			37196: outdata = 32'd28340;
			37197: outdata = 32'd28339;
			37198: outdata = 32'd28338;
			37199: outdata = 32'd28337;
			37200: outdata = 32'd28336;
			37201: outdata = 32'd28335;
			37202: outdata = 32'd28334;
			37203: outdata = 32'd28333;
			37204: outdata = 32'd28332;
			37205: outdata = 32'd28331;
			37206: outdata = 32'd28330;
			37207: outdata = 32'd28329;
			37208: outdata = 32'd28328;
			37209: outdata = 32'd28327;
			37210: outdata = 32'd28326;
			37211: outdata = 32'd28325;
			37212: outdata = 32'd28324;
			37213: outdata = 32'd28323;
			37214: outdata = 32'd28322;
			37215: outdata = 32'd28321;
			37216: outdata = 32'd28320;
			37217: outdata = 32'd28319;
			37218: outdata = 32'd28318;
			37219: outdata = 32'd28317;
			37220: outdata = 32'd28316;
			37221: outdata = 32'd28315;
			37222: outdata = 32'd28314;
			37223: outdata = 32'd28313;
			37224: outdata = 32'd28312;
			37225: outdata = 32'd28311;
			37226: outdata = 32'd28310;
			37227: outdata = 32'd28309;
			37228: outdata = 32'd28308;
			37229: outdata = 32'd28307;
			37230: outdata = 32'd28306;
			37231: outdata = 32'd28305;
			37232: outdata = 32'd28304;
			37233: outdata = 32'd28303;
			37234: outdata = 32'd28302;
			37235: outdata = 32'd28301;
			37236: outdata = 32'd28300;
			37237: outdata = 32'd28299;
			37238: outdata = 32'd28298;
			37239: outdata = 32'd28297;
			37240: outdata = 32'd28296;
			37241: outdata = 32'd28295;
			37242: outdata = 32'd28294;
			37243: outdata = 32'd28293;
			37244: outdata = 32'd28292;
			37245: outdata = 32'd28291;
			37246: outdata = 32'd28290;
			37247: outdata = 32'd28289;
			37248: outdata = 32'd28288;
			37249: outdata = 32'd28287;
			37250: outdata = 32'd28286;
			37251: outdata = 32'd28285;
			37252: outdata = 32'd28284;
			37253: outdata = 32'd28283;
			37254: outdata = 32'd28282;
			37255: outdata = 32'd28281;
			37256: outdata = 32'd28280;
			37257: outdata = 32'd28279;
			37258: outdata = 32'd28278;
			37259: outdata = 32'd28277;
			37260: outdata = 32'd28276;
			37261: outdata = 32'd28275;
			37262: outdata = 32'd28274;
			37263: outdata = 32'd28273;
			37264: outdata = 32'd28272;
			37265: outdata = 32'd28271;
			37266: outdata = 32'd28270;
			37267: outdata = 32'd28269;
			37268: outdata = 32'd28268;
			37269: outdata = 32'd28267;
			37270: outdata = 32'd28266;
			37271: outdata = 32'd28265;
			37272: outdata = 32'd28264;
			37273: outdata = 32'd28263;
			37274: outdata = 32'd28262;
			37275: outdata = 32'd28261;
			37276: outdata = 32'd28260;
			37277: outdata = 32'd28259;
			37278: outdata = 32'd28258;
			37279: outdata = 32'd28257;
			37280: outdata = 32'd28256;
			37281: outdata = 32'd28255;
			37282: outdata = 32'd28254;
			37283: outdata = 32'd28253;
			37284: outdata = 32'd28252;
			37285: outdata = 32'd28251;
			37286: outdata = 32'd28250;
			37287: outdata = 32'd28249;
			37288: outdata = 32'd28248;
			37289: outdata = 32'd28247;
			37290: outdata = 32'd28246;
			37291: outdata = 32'd28245;
			37292: outdata = 32'd28244;
			37293: outdata = 32'd28243;
			37294: outdata = 32'd28242;
			37295: outdata = 32'd28241;
			37296: outdata = 32'd28240;
			37297: outdata = 32'd28239;
			37298: outdata = 32'd28238;
			37299: outdata = 32'd28237;
			37300: outdata = 32'd28236;
			37301: outdata = 32'd28235;
			37302: outdata = 32'd28234;
			37303: outdata = 32'd28233;
			37304: outdata = 32'd28232;
			37305: outdata = 32'd28231;
			37306: outdata = 32'd28230;
			37307: outdata = 32'd28229;
			37308: outdata = 32'd28228;
			37309: outdata = 32'd28227;
			37310: outdata = 32'd28226;
			37311: outdata = 32'd28225;
			37312: outdata = 32'd28224;
			37313: outdata = 32'd28223;
			37314: outdata = 32'd28222;
			37315: outdata = 32'd28221;
			37316: outdata = 32'd28220;
			37317: outdata = 32'd28219;
			37318: outdata = 32'd28218;
			37319: outdata = 32'd28217;
			37320: outdata = 32'd28216;
			37321: outdata = 32'd28215;
			37322: outdata = 32'd28214;
			37323: outdata = 32'd28213;
			37324: outdata = 32'd28212;
			37325: outdata = 32'd28211;
			37326: outdata = 32'd28210;
			37327: outdata = 32'd28209;
			37328: outdata = 32'd28208;
			37329: outdata = 32'd28207;
			37330: outdata = 32'd28206;
			37331: outdata = 32'd28205;
			37332: outdata = 32'd28204;
			37333: outdata = 32'd28203;
			37334: outdata = 32'd28202;
			37335: outdata = 32'd28201;
			37336: outdata = 32'd28200;
			37337: outdata = 32'd28199;
			37338: outdata = 32'd28198;
			37339: outdata = 32'd28197;
			37340: outdata = 32'd28196;
			37341: outdata = 32'd28195;
			37342: outdata = 32'd28194;
			37343: outdata = 32'd28193;
			37344: outdata = 32'd28192;
			37345: outdata = 32'd28191;
			37346: outdata = 32'd28190;
			37347: outdata = 32'd28189;
			37348: outdata = 32'd28188;
			37349: outdata = 32'd28187;
			37350: outdata = 32'd28186;
			37351: outdata = 32'd28185;
			37352: outdata = 32'd28184;
			37353: outdata = 32'd28183;
			37354: outdata = 32'd28182;
			37355: outdata = 32'd28181;
			37356: outdata = 32'd28180;
			37357: outdata = 32'd28179;
			37358: outdata = 32'd28178;
			37359: outdata = 32'd28177;
			37360: outdata = 32'd28176;
			37361: outdata = 32'd28175;
			37362: outdata = 32'd28174;
			37363: outdata = 32'd28173;
			37364: outdata = 32'd28172;
			37365: outdata = 32'd28171;
			37366: outdata = 32'd28170;
			37367: outdata = 32'd28169;
			37368: outdata = 32'd28168;
			37369: outdata = 32'd28167;
			37370: outdata = 32'd28166;
			37371: outdata = 32'd28165;
			37372: outdata = 32'd28164;
			37373: outdata = 32'd28163;
			37374: outdata = 32'd28162;
			37375: outdata = 32'd28161;
			37376: outdata = 32'd28160;
			37377: outdata = 32'd28159;
			37378: outdata = 32'd28158;
			37379: outdata = 32'd28157;
			37380: outdata = 32'd28156;
			37381: outdata = 32'd28155;
			37382: outdata = 32'd28154;
			37383: outdata = 32'd28153;
			37384: outdata = 32'd28152;
			37385: outdata = 32'd28151;
			37386: outdata = 32'd28150;
			37387: outdata = 32'd28149;
			37388: outdata = 32'd28148;
			37389: outdata = 32'd28147;
			37390: outdata = 32'd28146;
			37391: outdata = 32'd28145;
			37392: outdata = 32'd28144;
			37393: outdata = 32'd28143;
			37394: outdata = 32'd28142;
			37395: outdata = 32'd28141;
			37396: outdata = 32'd28140;
			37397: outdata = 32'd28139;
			37398: outdata = 32'd28138;
			37399: outdata = 32'd28137;
			37400: outdata = 32'd28136;
			37401: outdata = 32'd28135;
			37402: outdata = 32'd28134;
			37403: outdata = 32'd28133;
			37404: outdata = 32'd28132;
			37405: outdata = 32'd28131;
			37406: outdata = 32'd28130;
			37407: outdata = 32'd28129;
			37408: outdata = 32'd28128;
			37409: outdata = 32'd28127;
			37410: outdata = 32'd28126;
			37411: outdata = 32'd28125;
			37412: outdata = 32'd28124;
			37413: outdata = 32'd28123;
			37414: outdata = 32'd28122;
			37415: outdata = 32'd28121;
			37416: outdata = 32'd28120;
			37417: outdata = 32'd28119;
			37418: outdata = 32'd28118;
			37419: outdata = 32'd28117;
			37420: outdata = 32'd28116;
			37421: outdata = 32'd28115;
			37422: outdata = 32'd28114;
			37423: outdata = 32'd28113;
			37424: outdata = 32'd28112;
			37425: outdata = 32'd28111;
			37426: outdata = 32'd28110;
			37427: outdata = 32'd28109;
			37428: outdata = 32'd28108;
			37429: outdata = 32'd28107;
			37430: outdata = 32'd28106;
			37431: outdata = 32'd28105;
			37432: outdata = 32'd28104;
			37433: outdata = 32'd28103;
			37434: outdata = 32'd28102;
			37435: outdata = 32'd28101;
			37436: outdata = 32'd28100;
			37437: outdata = 32'd28099;
			37438: outdata = 32'd28098;
			37439: outdata = 32'd28097;
			37440: outdata = 32'd28096;
			37441: outdata = 32'd28095;
			37442: outdata = 32'd28094;
			37443: outdata = 32'd28093;
			37444: outdata = 32'd28092;
			37445: outdata = 32'd28091;
			37446: outdata = 32'd28090;
			37447: outdata = 32'd28089;
			37448: outdata = 32'd28088;
			37449: outdata = 32'd28087;
			37450: outdata = 32'd28086;
			37451: outdata = 32'd28085;
			37452: outdata = 32'd28084;
			37453: outdata = 32'd28083;
			37454: outdata = 32'd28082;
			37455: outdata = 32'd28081;
			37456: outdata = 32'd28080;
			37457: outdata = 32'd28079;
			37458: outdata = 32'd28078;
			37459: outdata = 32'd28077;
			37460: outdata = 32'd28076;
			37461: outdata = 32'd28075;
			37462: outdata = 32'd28074;
			37463: outdata = 32'd28073;
			37464: outdata = 32'd28072;
			37465: outdata = 32'd28071;
			37466: outdata = 32'd28070;
			37467: outdata = 32'd28069;
			37468: outdata = 32'd28068;
			37469: outdata = 32'd28067;
			37470: outdata = 32'd28066;
			37471: outdata = 32'd28065;
			37472: outdata = 32'd28064;
			37473: outdata = 32'd28063;
			37474: outdata = 32'd28062;
			37475: outdata = 32'd28061;
			37476: outdata = 32'd28060;
			37477: outdata = 32'd28059;
			37478: outdata = 32'd28058;
			37479: outdata = 32'd28057;
			37480: outdata = 32'd28056;
			37481: outdata = 32'd28055;
			37482: outdata = 32'd28054;
			37483: outdata = 32'd28053;
			37484: outdata = 32'd28052;
			37485: outdata = 32'd28051;
			37486: outdata = 32'd28050;
			37487: outdata = 32'd28049;
			37488: outdata = 32'd28048;
			37489: outdata = 32'd28047;
			37490: outdata = 32'd28046;
			37491: outdata = 32'd28045;
			37492: outdata = 32'd28044;
			37493: outdata = 32'd28043;
			37494: outdata = 32'd28042;
			37495: outdata = 32'd28041;
			37496: outdata = 32'd28040;
			37497: outdata = 32'd28039;
			37498: outdata = 32'd28038;
			37499: outdata = 32'd28037;
			37500: outdata = 32'd28036;
			37501: outdata = 32'd28035;
			37502: outdata = 32'd28034;
			37503: outdata = 32'd28033;
			37504: outdata = 32'd28032;
			37505: outdata = 32'd28031;
			37506: outdata = 32'd28030;
			37507: outdata = 32'd28029;
			37508: outdata = 32'd28028;
			37509: outdata = 32'd28027;
			37510: outdata = 32'd28026;
			37511: outdata = 32'd28025;
			37512: outdata = 32'd28024;
			37513: outdata = 32'd28023;
			37514: outdata = 32'd28022;
			37515: outdata = 32'd28021;
			37516: outdata = 32'd28020;
			37517: outdata = 32'd28019;
			37518: outdata = 32'd28018;
			37519: outdata = 32'd28017;
			37520: outdata = 32'd28016;
			37521: outdata = 32'd28015;
			37522: outdata = 32'd28014;
			37523: outdata = 32'd28013;
			37524: outdata = 32'd28012;
			37525: outdata = 32'd28011;
			37526: outdata = 32'd28010;
			37527: outdata = 32'd28009;
			37528: outdata = 32'd28008;
			37529: outdata = 32'd28007;
			37530: outdata = 32'd28006;
			37531: outdata = 32'd28005;
			37532: outdata = 32'd28004;
			37533: outdata = 32'd28003;
			37534: outdata = 32'd28002;
			37535: outdata = 32'd28001;
			37536: outdata = 32'd28000;
			37537: outdata = 32'd27999;
			37538: outdata = 32'd27998;
			37539: outdata = 32'd27997;
			37540: outdata = 32'd27996;
			37541: outdata = 32'd27995;
			37542: outdata = 32'd27994;
			37543: outdata = 32'd27993;
			37544: outdata = 32'd27992;
			37545: outdata = 32'd27991;
			37546: outdata = 32'd27990;
			37547: outdata = 32'd27989;
			37548: outdata = 32'd27988;
			37549: outdata = 32'd27987;
			37550: outdata = 32'd27986;
			37551: outdata = 32'd27985;
			37552: outdata = 32'd27984;
			37553: outdata = 32'd27983;
			37554: outdata = 32'd27982;
			37555: outdata = 32'd27981;
			37556: outdata = 32'd27980;
			37557: outdata = 32'd27979;
			37558: outdata = 32'd27978;
			37559: outdata = 32'd27977;
			37560: outdata = 32'd27976;
			37561: outdata = 32'd27975;
			37562: outdata = 32'd27974;
			37563: outdata = 32'd27973;
			37564: outdata = 32'd27972;
			37565: outdata = 32'd27971;
			37566: outdata = 32'd27970;
			37567: outdata = 32'd27969;
			37568: outdata = 32'd27968;
			37569: outdata = 32'd27967;
			37570: outdata = 32'd27966;
			37571: outdata = 32'd27965;
			37572: outdata = 32'd27964;
			37573: outdata = 32'd27963;
			37574: outdata = 32'd27962;
			37575: outdata = 32'd27961;
			37576: outdata = 32'd27960;
			37577: outdata = 32'd27959;
			37578: outdata = 32'd27958;
			37579: outdata = 32'd27957;
			37580: outdata = 32'd27956;
			37581: outdata = 32'd27955;
			37582: outdata = 32'd27954;
			37583: outdata = 32'd27953;
			37584: outdata = 32'd27952;
			37585: outdata = 32'd27951;
			37586: outdata = 32'd27950;
			37587: outdata = 32'd27949;
			37588: outdata = 32'd27948;
			37589: outdata = 32'd27947;
			37590: outdata = 32'd27946;
			37591: outdata = 32'd27945;
			37592: outdata = 32'd27944;
			37593: outdata = 32'd27943;
			37594: outdata = 32'd27942;
			37595: outdata = 32'd27941;
			37596: outdata = 32'd27940;
			37597: outdata = 32'd27939;
			37598: outdata = 32'd27938;
			37599: outdata = 32'd27937;
			37600: outdata = 32'd27936;
			37601: outdata = 32'd27935;
			37602: outdata = 32'd27934;
			37603: outdata = 32'd27933;
			37604: outdata = 32'd27932;
			37605: outdata = 32'd27931;
			37606: outdata = 32'd27930;
			37607: outdata = 32'd27929;
			37608: outdata = 32'd27928;
			37609: outdata = 32'd27927;
			37610: outdata = 32'd27926;
			37611: outdata = 32'd27925;
			37612: outdata = 32'd27924;
			37613: outdata = 32'd27923;
			37614: outdata = 32'd27922;
			37615: outdata = 32'd27921;
			37616: outdata = 32'd27920;
			37617: outdata = 32'd27919;
			37618: outdata = 32'd27918;
			37619: outdata = 32'd27917;
			37620: outdata = 32'd27916;
			37621: outdata = 32'd27915;
			37622: outdata = 32'd27914;
			37623: outdata = 32'd27913;
			37624: outdata = 32'd27912;
			37625: outdata = 32'd27911;
			37626: outdata = 32'd27910;
			37627: outdata = 32'd27909;
			37628: outdata = 32'd27908;
			37629: outdata = 32'd27907;
			37630: outdata = 32'd27906;
			37631: outdata = 32'd27905;
			37632: outdata = 32'd27904;
			37633: outdata = 32'd27903;
			37634: outdata = 32'd27902;
			37635: outdata = 32'd27901;
			37636: outdata = 32'd27900;
			37637: outdata = 32'd27899;
			37638: outdata = 32'd27898;
			37639: outdata = 32'd27897;
			37640: outdata = 32'd27896;
			37641: outdata = 32'd27895;
			37642: outdata = 32'd27894;
			37643: outdata = 32'd27893;
			37644: outdata = 32'd27892;
			37645: outdata = 32'd27891;
			37646: outdata = 32'd27890;
			37647: outdata = 32'd27889;
			37648: outdata = 32'd27888;
			37649: outdata = 32'd27887;
			37650: outdata = 32'd27886;
			37651: outdata = 32'd27885;
			37652: outdata = 32'd27884;
			37653: outdata = 32'd27883;
			37654: outdata = 32'd27882;
			37655: outdata = 32'd27881;
			37656: outdata = 32'd27880;
			37657: outdata = 32'd27879;
			37658: outdata = 32'd27878;
			37659: outdata = 32'd27877;
			37660: outdata = 32'd27876;
			37661: outdata = 32'd27875;
			37662: outdata = 32'd27874;
			37663: outdata = 32'd27873;
			37664: outdata = 32'd27872;
			37665: outdata = 32'd27871;
			37666: outdata = 32'd27870;
			37667: outdata = 32'd27869;
			37668: outdata = 32'd27868;
			37669: outdata = 32'd27867;
			37670: outdata = 32'd27866;
			37671: outdata = 32'd27865;
			37672: outdata = 32'd27864;
			37673: outdata = 32'd27863;
			37674: outdata = 32'd27862;
			37675: outdata = 32'd27861;
			37676: outdata = 32'd27860;
			37677: outdata = 32'd27859;
			37678: outdata = 32'd27858;
			37679: outdata = 32'd27857;
			37680: outdata = 32'd27856;
			37681: outdata = 32'd27855;
			37682: outdata = 32'd27854;
			37683: outdata = 32'd27853;
			37684: outdata = 32'd27852;
			37685: outdata = 32'd27851;
			37686: outdata = 32'd27850;
			37687: outdata = 32'd27849;
			37688: outdata = 32'd27848;
			37689: outdata = 32'd27847;
			37690: outdata = 32'd27846;
			37691: outdata = 32'd27845;
			37692: outdata = 32'd27844;
			37693: outdata = 32'd27843;
			37694: outdata = 32'd27842;
			37695: outdata = 32'd27841;
			37696: outdata = 32'd27840;
			37697: outdata = 32'd27839;
			37698: outdata = 32'd27838;
			37699: outdata = 32'd27837;
			37700: outdata = 32'd27836;
			37701: outdata = 32'd27835;
			37702: outdata = 32'd27834;
			37703: outdata = 32'd27833;
			37704: outdata = 32'd27832;
			37705: outdata = 32'd27831;
			37706: outdata = 32'd27830;
			37707: outdata = 32'd27829;
			37708: outdata = 32'd27828;
			37709: outdata = 32'd27827;
			37710: outdata = 32'd27826;
			37711: outdata = 32'd27825;
			37712: outdata = 32'd27824;
			37713: outdata = 32'd27823;
			37714: outdata = 32'd27822;
			37715: outdata = 32'd27821;
			37716: outdata = 32'd27820;
			37717: outdata = 32'd27819;
			37718: outdata = 32'd27818;
			37719: outdata = 32'd27817;
			37720: outdata = 32'd27816;
			37721: outdata = 32'd27815;
			37722: outdata = 32'd27814;
			37723: outdata = 32'd27813;
			37724: outdata = 32'd27812;
			37725: outdata = 32'd27811;
			37726: outdata = 32'd27810;
			37727: outdata = 32'd27809;
			37728: outdata = 32'd27808;
			37729: outdata = 32'd27807;
			37730: outdata = 32'd27806;
			37731: outdata = 32'd27805;
			37732: outdata = 32'd27804;
			37733: outdata = 32'd27803;
			37734: outdata = 32'd27802;
			37735: outdata = 32'd27801;
			37736: outdata = 32'd27800;
			37737: outdata = 32'd27799;
			37738: outdata = 32'd27798;
			37739: outdata = 32'd27797;
			37740: outdata = 32'd27796;
			37741: outdata = 32'd27795;
			37742: outdata = 32'd27794;
			37743: outdata = 32'd27793;
			37744: outdata = 32'd27792;
			37745: outdata = 32'd27791;
			37746: outdata = 32'd27790;
			37747: outdata = 32'd27789;
			37748: outdata = 32'd27788;
			37749: outdata = 32'd27787;
			37750: outdata = 32'd27786;
			37751: outdata = 32'd27785;
			37752: outdata = 32'd27784;
			37753: outdata = 32'd27783;
			37754: outdata = 32'd27782;
			37755: outdata = 32'd27781;
			37756: outdata = 32'd27780;
			37757: outdata = 32'd27779;
			37758: outdata = 32'd27778;
			37759: outdata = 32'd27777;
			37760: outdata = 32'd27776;
			37761: outdata = 32'd27775;
			37762: outdata = 32'd27774;
			37763: outdata = 32'd27773;
			37764: outdata = 32'd27772;
			37765: outdata = 32'd27771;
			37766: outdata = 32'd27770;
			37767: outdata = 32'd27769;
			37768: outdata = 32'd27768;
			37769: outdata = 32'd27767;
			37770: outdata = 32'd27766;
			37771: outdata = 32'd27765;
			37772: outdata = 32'd27764;
			37773: outdata = 32'd27763;
			37774: outdata = 32'd27762;
			37775: outdata = 32'd27761;
			37776: outdata = 32'd27760;
			37777: outdata = 32'd27759;
			37778: outdata = 32'd27758;
			37779: outdata = 32'd27757;
			37780: outdata = 32'd27756;
			37781: outdata = 32'd27755;
			37782: outdata = 32'd27754;
			37783: outdata = 32'd27753;
			37784: outdata = 32'd27752;
			37785: outdata = 32'd27751;
			37786: outdata = 32'd27750;
			37787: outdata = 32'd27749;
			37788: outdata = 32'd27748;
			37789: outdata = 32'd27747;
			37790: outdata = 32'd27746;
			37791: outdata = 32'd27745;
			37792: outdata = 32'd27744;
			37793: outdata = 32'd27743;
			37794: outdata = 32'd27742;
			37795: outdata = 32'd27741;
			37796: outdata = 32'd27740;
			37797: outdata = 32'd27739;
			37798: outdata = 32'd27738;
			37799: outdata = 32'd27737;
			37800: outdata = 32'd27736;
			37801: outdata = 32'd27735;
			37802: outdata = 32'd27734;
			37803: outdata = 32'd27733;
			37804: outdata = 32'd27732;
			37805: outdata = 32'd27731;
			37806: outdata = 32'd27730;
			37807: outdata = 32'd27729;
			37808: outdata = 32'd27728;
			37809: outdata = 32'd27727;
			37810: outdata = 32'd27726;
			37811: outdata = 32'd27725;
			37812: outdata = 32'd27724;
			37813: outdata = 32'd27723;
			37814: outdata = 32'd27722;
			37815: outdata = 32'd27721;
			37816: outdata = 32'd27720;
			37817: outdata = 32'd27719;
			37818: outdata = 32'd27718;
			37819: outdata = 32'd27717;
			37820: outdata = 32'd27716;
			37821: outdata = 32'd27715;
			37822: outdata = 32'd27714;
			37823: outdata = 32'd27713;
			37824: outdata = 32'd27712;
			37825: outdata = 32'd27711;
			37826: outdata = 32'd27710;
			37827: outdata = 32'd27709;
			37828: outdata = 32'd27708;
			37829: outdata = 32'd27707;
			37830: outdata = 32'd27706;
			37831: outdata = 32'd27705;
			37832: outdata = 32'd27704;
			37833: outdata = 32'd27703;
			37834: outdata = 32'd27702;
			37835: outdata = 32'd27701;
			37836: outdata = 32'd27700;
			37837: outdata = 32'd27699;
			37838: outdata = 32'd27698;
			37839: outdata = 32'd27697;
			37840: outdata = 32'd27696;
			37841: outdata = 32'd27695;
			37842: outdata = 32'd27694;
			37843: outdata = 32'd27693;
			37844: outdata = 32'd27692;
			37845: outdata = 32'd27691;
			37846: outdata = 32'd27690;
			37847: outdata = 32'd27689;
			37848: outdata = 32'd27688;
			37849: outdata = 32'd27687;
			37850: outdata = 32'd27686;
			37851: outdata = 32'd27685;
			37852: outdata = 32'd27684;
			37853: outdata = 32'd27683;
			37854: outdata = 32'd27682;
			37855: outdata = 32'd27681;
			37856: outdata = 32'd27680;
			37857: outdata = 32'd27679;
			37858: outdata = 32'd27678;
			37859: outdata = 32'd27677;
			37860: outdata = 32'd27676;
			37861: outdata = 32'd27675;
			37862: outdata = 32'd27674;
			37863: outdata = 32'd27673;
			37864: outdata = 32'd27672;
			37865: outdata = 32'd27671;
			37866: outdata = 32'd27670;
			37867: outdata = 32'd27669;
			37868: outdata = 32'd27668;
			37869: outdata = 32'd27667;
			37870: outdata = 32'd27666;
			37871: outdata = 32'd27665;
			37872: outdata = 32'd27664;
			37873: outdata = 32'd27663;
			37874: outdata = 32'd27662;
			37875: outdata = 32'd27661;
			37876: outdata = 32'd27660;
			37877: outdata = 32'd27659;
			37878: outdata = 32'd27658;
			37879: outdata = 32'd27657;
			37880: outdata = 32'd27656;
			37881: outdata = 32'd27655;
			37882: outdata = 32'd27654;
			37883: outdata = 32'd27653;
			37884: outdata = 32'd27652;
			37885: outdata = 32'd27651;
			37886: outdata = 32'd27650;
			37887: outdata = 32'd27649;
			37888: outdata = 32'd27648;
			37889: outdata = 32'd27647;
			37890: outdata = 32'd27646;
			37891: outdata = 32'd27645;
			37892: outdata = 32'd27644;
			37893: outdata = 32'd27643;
			37894: outdata = 32'd27642;
			37895: outdata = 32'd27641;
			37896: outdata = 32'd27640;
			37897: outdata = 32'd27639;
			37898: outdata = 32'd27638;
			37899: outdata = 32'd27637;
			37900: outdata = 32'd27636;
			37901: outdata = 32'd27635;
			37902: outdata = 32'd27634;
			37903: outdata = 32'd27633;
			37904: outdata = 32'd27632;
			37905: outdata = 32'd27631;
			37906: outdata = 32'd27630;
			37907: outdata = 32'd27629;
			37908: outdata = 32'd27628;
			37909: outdata = 32'd27627;
			37910: outdata = 32'd27626;
			37911: outdata = 32'd27625;
			37912: outdata = 32'd27624;
			37913: outdata = 32'd27623;
			37914: outdata = 32'd27622;
			37915: outdata = 32'd27621;
			37916: outdata = 32'd27620;
			37917: outdata = 32'd27619;
			37918: outdata = 32'd27618;
			37919: outdata = 32'd27617;
			37920: outdata = 32'd27616;
			37921: outdata = 32'd27615;
			37922: outdata = 32'd27614;
			37923: outdata = 32'd27613;
			37924: outdata = 32'd27612;
			37925: outdata = 32'd27611;
			37926: outdata = 32'd27610;
			37927: outdata = 32'd27609;
			37928: outdata = 32'd27608;
			37929: outdata = 32'd27607;
			37930: outdata = 32'd27606;
			37931: outdata = 32'd27605;
			37932: outdata = 32'd27604;
			37933: outdata = 32'd27603;
			37934: outdata = 32'd27602;
			37935: outdata = 32'd27601;
			37936: outdata = 32'd27600;
			37937: outdata = 32'd27599;
			37938: outdata = 32'd27598;
			37939: outdata = 32'd27597;
			37940: outdata = 32'd27596;
			37941: outdata = 32'd27595;
			37942: outdata = 32'd27594;
			37943: outdata = 32'd27593;
			37944: outdata = 32'd27592;
			37945: outdata = 32'd27591;
			37946: outdata = 32'd27590;
			37947: outdata = 32'd27589;
			37948: outdata = 32'd27588;
			37949: outdata = 32'd27587;
			37950: outdata = 32'd27586;
			37951: outdata = 32'd27585;
			37952: outdata = 32'd27584;
			37953: outdata = 32'd27583;
			37954: outdata = 32'd27582;
			37955: outdata = 32'd27581;
			37956: outdata = 32'd27580;
			37957: outdata = 32'd27579;
			37958: outdata = 32'd27578;
			37959: outdata = 32'd27577;
			37960: outdata = 32'd27576;
			37961: outdata = 32'd27575;
			37962: outdata = 32'd27574;
			37963: outdata = 32'd27573;
			37964: outdata = 32'd27572;
			37965: outdata = 32'd27571;
			37966: outdata = 32'd27570;
			37967: outdata = 32'd27569;
			37968: outdata = 32'd27568;
			37969: outdata = 32'd27567;
			37970: outdata = 32'd27566;
			37971: outdata = 32'd27565;
			37972: outdata = 32'd27564;
			37973: outdata = 32'd27563;
			37974: outdata = 32'd27562;
			37975: outdata = 32'd27561;
			37976: outdata = 32'd27560;
			37977: outdata = 32'd27559;
			37978: outdata = 32'd27558;
			37979: outdata = 32'd27557;
			37980: outdata = 32'd27556;
			37981: outdata = 32'd27555;
			37982: outdata = 32'd27554;
			37983: outdata = 32'd27553;
			37984: outdata = 32'd27552;
			37985: outdata = 32'd27551;
			37986: outdata = 32'd27550;
			37987: outdata = 32'd27549;
			37988: outdata = 32'd27548;
			37989: outdata = 32'd27547;
			37990: outdata = 32'd27546;
			37991: outdata = 32'd27545;
			37992: outdata = 32'd27544;
			37993: outdata = 32'd27543;
			37994: outdata = 32'd27542;
			37995: outdata = 32'd27541;
			37996: outdata = 32'd27540;
			37997: outdata = 32'd27539;
			37998: outdata = 32'd27538;
			37999: outdata = 32'd27537;
			38000: outdata = 32'd27536;
			38001: outdata = 32'd27535;
			38002: outdata = 32'd27534;
			38003: outdata = 32'd27533;
			38004: outdata = 32'd27532;
			38005: outdata = 32'd27531;
			38006: outdata = 32'd27530;
			38007: outdata = 32'd27529;
			38008: outdata = 32'd27528;
			38009: outdata = 32'd27527;
			38010: outdata = 32'd27526;
			38011: outdata = 32'd27525;
			38012: outdata = 32'd27524;
			38013: outdata = 32'd27523;
			38014: outdata = 32'd27522;
			38015: outdata = 32'd27521;
			38016: outdata = 32'd27520;
			38017: outdata = 32'd27519;
			38018: outdata = 32'd27518;
			38019: outdata = 32'd27517;
			38020: outdata = 32'd27516;
			38021: outdata = 32'd27515;
			38022: outdata = 32'd27514;
			38023: outdata = 32'd27513;
			38024: outdata = 32'd27512;
			38025: outdata = 32'd27511;
			38026: outdata = 32'd27510;
			38027: outdata = 32'd27509;
			38028: outdata = 32'd27508;
			38029: outdata = 32'd27507;
			38030: outdata = 32'd27506;
			38031: outdata = 32'd27505;
			38032: outdata = 32'd27504;
			38033: outdata = 32'd27503;
			38034: outdata = 32'd27502;
			38035: outdata = 32'd27501;
			38036: outdata = 32'd27500;
			38037: outdata = 32'd27499;
			38038: outdata = 32'd27498;
			38039: outdata = 32'd27497;
			38040: outdata = 32'd27496;
			38041: outdata = 32'd27495;
			38042: outdata = 32'd27494;
			38043: outdata = 32'd27493;
			38044: outdata = 32'd27492;
			38045: outdata = 32'd27491;
			38046: outdata = 32'd27490;
			38047: outdata = 32'd27489;
			38048: outdata = 32'd27488;
			38049: outdata = 32'd27487;
			38050: outdata = 32'd27486;
			38051: outdata = 32'd27485;
			38052: outdata = 32'd27484;
			38053: outdata = 32'd27483;
			38054: outdata = 32'd27482;
			38055: outdata = 32'd27481;
			38056: outdata = 32'd27480;
			38057: outdata = 32'd27479;
			38058: outdata = 32'd27478;
			38059: outdata = 32'd27477;
			38060: outdata = 32'd27476;
			38061: outdata = 32'd27475;
			38062: outdata = 32'd27474;
			38063: outdata = 32'd27473;
			38064: outdata = 32'd27472;
			38065: outdata = 32'd27471;
			38066: outdata = 32'd27470;
			38067: outdata = 32'd27469;
			38068: outdata = 32'd27468;
			38069: outdata = 32'd27467;
			38070: outdata = 32'd27466;
			38071: outdata = 32'd27465;
			38072: outdata = 32'd27464;
			38073: outdata = 32'd27463;
			38074: outdata = 32'd27462;
			38075: outdata = 32'd27461;
			38076: outdata = 32'd27460;
			38077: outdata = 32'd27459;
			38078: outdata = 32'd27458;
			38079: outdata = 32'd27457;
			38080: outdata = 32'd27456;
			38081: outdata = 32'd27455;
			38082: outdata = 32'd27454;
			38083: outdata = 32'd27453;
			38084: outdata = 32'd27452;
			38085: outdata = 32'd27451;
			38086: outdata = 32'd27450;
			38087: outdata = 32'd27449;
			38088: outdata = 32'd27448;
			38089: outdata = 32'd27447;
			38090: outdata = 32'd27446;
			38091: outdata = 32'd27445;
			38092: outdata = 32'd27444;
			38093: outdata = 32'd27443;
			38094: outdata = 32'd27442;
			38095: outdata = 32'd27441;
			38096: outdata = 32'd27440;
			38097: outdata = 32'd27439;
			38098: outdata = 32'd27438;
			38099: outdata = 32'd27437;
			38100: outdata = 32'd27436;
			38101: outdata = 32'd27435;
			38102: outdata = 32'd27434;
			38103: outdata = 32'd27433;
			38104: outdata = 32'd27432;
			38105: outdata = 32'd27431;
			38106: outdata = 32'd27430;
			38107: outdata = 32'd27429;
			38108: outdata = 32'd27428;
			38109: outdata = 32'd27427;
			38110: outdata = 32'd27426;
			38111: outdata = 32'd27425;
			38112: outdata = 32'd27424;
			38113: outdata = 32'd27423;
			38114: outdata = 32'd27422;
			38115: outdata = 32'd27421;
			38116: outdata = 32'd27420;
			38117: outdata = 32'd27419;
			38118: outdata = 32'd27418;
			38119: outdata = 32'd27417;
			38120: outdata = 32'd27416;
			38121: outdata = 32'd27415;
			38122: outdata = 32'd27414;
			38123: outdata = 32'd27413;
			38124: outdata = 32'd27412;
			38125: outdata = 32'd27411;
			38126: outdata = 32'd27410;
			38127: outdata = 32'd27409;
			38128: outdata = 32'd27408;
			38129: outdata = 32'd27407;
			38130: outdata = 32'd27406;
			38131: outdata = 32'd27405;
			38132: outdata = 32'd27404;
			38133: outdata = 32'd27403;
			38134: outdata = 32'd27402;
			38135: outdata = 32'd27401;
			38136: outdata = 32'd27400;
			38137: outdata = 32'd27399;
			38138: outdata = 32'd27398;
			38139: outdata = 32'd27397;
			38140: outdata = 32'd27396;
			38141: outdata = 32'd27395;
			38142: outdata = 32'd27394;
			38143: outdata = 32'd27393;
			38144: outdata = 32'd27392;
			38145: outdata = 32'd27391;
			38146: outdata = 32'd27390;
			38147: outdata = 32'd27389;
			38148: outdata = 32'd27388;
			38149: outdata = 32'd27387;
			38150: outdata = 32'd27386;
			38151: outdata = 32'd27385;
			38152: outdata = 32'd27384;
			38153: outdata = 32'd27383;
			38154: outdata = 32'd27382;
			38155: outdata = 32'd27381;
			38156: outdata = 32'd27380;
			38157: outdata = 32'd27379;
			38158: outdata = 32'd27378;
			38159: outdata = 32'd27377;
			38160: outdata = 32'd27376;
			38161: outdata = 32'd27375;
			38162: outdata = 32'd27374;
			38163: outdata = 32'd27373;
			38164: outdata = 32'd27372;
			38165: outdata = 32'd27371;
			38166: outdata = 32'd27370;
			38167: outdata = 32'd27369;
			38168: outdata = 32'd27368;
			38169: outdata = 32'd27367;
			38170: outdata = 32'd27366;
			38171: outdata = 32'd27365;
			38172: outdata = 32'd27364;
			38173: outdata = 32'd27363;
			38174: outdata = 32'd27362;
			38175: outdata = 32'd27361;
			38176: outdata = 32'd27360;
			38177: outdata = 32'd27359;
			38178: outdata = 32'd27358;
			38179: outdata = 32'd27357;
			38180: outdata = 32'd27356;
			38181: outdata = 32'd27355;
			38182: outdata = 32'd27354;
			38183: outdata = 32'd27353;
			38184: outdata = 32'd27352;
			38185: outdata = 32'd27351;
			38186: outdata = 32'd27350;
			38187: outdata = 32'd27349;
			38188: outdata = 32'd27348;
			38189: outdata = 32'd27347;
			38190: outdata = 32'd27346;
			38191: outdata = 32'd27345;
			38192: outdata = 32'd27344;
			38193: outdata = 32'd27343;
			38194: outdata = 32'd27342;
			38195: outdata = 32'd27341;
			38196: outdata = 32'd27340;
			38197: outdata = 32'd27339;
			38198: outdata = 32'd27338;
			38199: outdata = 32'd27337;
			38200: outdata = 32'd27336;
			38201: outdata = 32'd27335;
			38202: outdata = 32'd27334;
			38203: outdata = 32'd27333;
			38204: outdata = 32'd27332;
			38205: outdata = 32'd27331;
			38206: outdata = 32'd27330;
			38207: outdata = 32'd27329;
			38208: outdata = 32'd27328;
			38209: outdata = 32'd27327;
			38210: outdata = 32'd27326;
			38211: outdata = 32'd27325;
			38212: outdata = 32'd27324;
			38213: outdata = 32'd27323;
			38214: outdata = 32'd27322;
			38215: outdata = 32'd27321;
			38216: outdata = 32'd27320;
			38217: outdata = 32'd27319;
			38218: outdata = 32'd27318;
			38219: outdata = 32'd27317;
			38220: outdata = 32'd27316;
			38221: outdata = 32'd27315;
			38222: outdata = 32'd27314;
			38223: outdata = 32'd27313;
			38224: outdata = 32'd27312;
			38225: outdata = 32'd27311;
			38226: outdata = 32'd27310;
			38227: outdata = 32'd27309;
			38228: outdata = 32'd27308;
			38229: outdata = 32'd27307;
			38230: outdata = 32'd27306;
			38231: outdata = 32'd27305;
			38232: outdata = 32'd27304;
			38233: outdata = 32'd27303;
			38234: outdata = 32'd27302;
			38235: outdata = 32'd27301;
			38236: outdata = 32'd27300;
			38237: outdata = 32'd27299;
			38238: outdata = 32'd27298;
			38239: outdata = 32'd27297;
			38240: outdata = 32'd27296;
			38241: outdata = 32'd27295;
			38242: outdata = 32'd27294;
			38243: outdata = 32'd27293;
			38244: outdata = 32'd27292;
			38245: outdata = 32'd27291;
			38246: outdata = 32'd27290;
			38247: outdata = 32'd27289;
			38248: outdata = 32'd27288;
			38249: outdata = 32'd27287;
			38250: outdata = 32'd27286;
			38251: outdata = 32'd27285;
			38252: outdata = 32'd27284;
			38253: outdata = 32'd27283;
			38254: outdata = 32'd27282;
			38255: outdata = 32'd27281;
			38256: outdata = 32'd27280;
			38257: outdata = 32'd27279;
			38258: outdata = 32'd27278;
			38259: outdata = 32'd27277;
			38260: outdata = 32'd27276;
			38261: outdata = 32'd27275;
			38262: outdata = 32'd27274;
			38263: outdata = 32'd27273;
			38264: outdata = 32'd27272;
			38265: outdata = 32'd27271;
			38266: outdata = 32'd27270;
			38267: outdata = 32'd27269;
			38268: outdata = 32'd27268;
			38269: outdata = 32'd27267;
			38270: outdata = 32'd27266;
			38271: outdata = 32'd27265;
			38272: outdata = 32'd27264;
			38273: outdata = 32'd27263;
			38274: outdata = 32'd27262;
			38275: outdata = 32'd27261;
			38276: outdata = 32'd27260;
			38277: outdata = 32'd27259;
			38278: outdata = 32'd27258;
			38279: outdata = 32'd27257;
			38280: outdata = 32'd27256;
			38281: outdata = 32'd27255;
			38282: outdata = 32'd27254;
			38283: outdata = 32'd27253;
			38284: outdata = 32'd27252;
			38285: outdata = 32'd27251;
			38286: outdata = 32'd27250;
			38287: outdata = 32'd27249;
			38288: outdata = 32'd27248;
			38289: outdata = 32'd27247;
			38290: outdata = 32'd27246;
			38291: outdata = 32'd27245;
			38292: outdata = 32'd27244;
			38293: outdata = 32'd27243;
			38294: outdata = 32'd27242;
			38295: outdata = 32'd27241;
			38296: outdata = 32'd27240;
			38297: outdata = 32'd27239;
			38298: outdata = 32'd27238;
			38299: outdata = 32'd27237;
			38300: outdata = 32'd27236;
			38301: outdata = 32'd27235;
			38302: outdata = 32'd27234;
			38303: outdata = 32'd27233;
			38304: outdata = 32'd27232;
			38305: outdata = 32'd27231;
			38306: outdata = 32'd27230;
			38307: outdata = 32'd27229;
			38308: outdata = 32'd27228;
			38309: outdata = 32'd27227;
			38310: outdata = 32'd27226;
			38311: outdata = 32'd27225;
			38312: outdata = 32'd27224;
			38313: outdata = 32'd27223;
			38314: outdata = 32'd27222;
			38315: outdata = 32'd27221;
			38316: outdata = 32'd27220;
			38317: outdata = 32'd27219;
			38318: outdata = 32'd27218;
			38319: outdata = 32'd27217;
			38320: outdata = 32'd27216;
			38321: outdata = 32'd27215;
			38322: outdata = 32'd27214;
			38323: outdata = 32'd27213;
			38324: outdata = 32'd27212;
			38325: outdata = 32'd27211;
			38326: outdata = 32'd27210;
			38327: outdata = 32'd27209;
			38328: outdata = 32'd27208;
			38329: outdata = 32'd27207;
			38330: outdata = 32'd27206;
			38331: outdata = 32'd27205;
			38332: outdata = 32'd27204;
			38333: outdata = 32'd27203;
			38334: outdata = 32'd27202;
			38335: outdata = 32'd27201;
			38336: outdata = 32'd27200;
			38337: outdata = 32'd27199;
			38338: outdata = 32'd27198;
			38339: outdata = 32'd27197;
			38340: outdata = 32'd27196;
			38341: outdata = 32'd27195;
			38342: outdata = 32'd27194;
			38343: outdata = 32'd27193;
			38344: outdata = 32'd27192;
			38345: outdata = 32'd27191;
			38346: outdata = 32'd27190;
			38347: outdata = 32'd27189;
			38348: outdata = 32'd27188;
			38349: outdata = 32'd27187;
			38350: outdata = 32'd27186;
			38351: outdata = 32'd27185;
			38352: outdata = 32'd27184;
			38353: outdata = 32'd27183;
			38354: outdata = 32'd27182;
			38355: outdata = 32'd27181;
			38356: outdata = 32'd27180;
			38357: outdata = 32'd27179;
			38358: outdata = 32'd27178;
			38359: outdata = 32'd27177;
			38360: outdata = 32'd27176;
			38361: outdata = 32'd27175;
			38362: outdata = 32'd27174;
			38363: outdata = 32'd27173;
			38364: outdata = 32'd27172;
			38365: outdata = 32'd27171;
			38366: outdata = 32'd27170;
			38367: outdata = 32'd27169;
			38368: outdata = 32'd27168;
			38369: outdata = 32'd27167;
			38370: outdata = 32'd27166;
			38371: outdata = 32'd27165;
			38372: outdata = 32'd27164;
			38373: outdata = 32'd27163;
			38374: outdata = 32'd27162;
			38375: outdata = 32'd27161;
			38376: outdata = 32'd27160;
			38377: outdata = 32'd27159;
			38378: outdata = 32'd27158;
			38379: outdata = 32'd27157;
			38380: outdata = 32'd27156;
			38381: outdata = 32'd27155;
			38382: outdata = 32'd27154;
			38383: outdata = 32'd27153;
			38384: outdata = 32'd27152;
			38385: outdata = 32'd27151;
			38386: outdata = 32'd27150;
			38387: outdata = 32'd27149;
			38388: outdata = 32'd27148;
			38389: outdata = 32'd27147;
			38390: outdata = 32'd27146;
			38391: outdata = 32'd27145;
			38392: outdata = 32'd27144;
			38393: outdata = 32'd27143;
			38394: outdata = 32'd27142;
			38395: outdata = 32'd27141;
			38396: outdata = 32'd27140;
			38397: outdata = 32'd27139;
			38398: outdata = 32'd27138;
			38399: outdata = 32'd27137;
			38400: outdata = 32'd27136;
			38401: outdata = 32'd27135;
			38402: outdata = 32'd27134;
			38403: outdata = 32'd27133;
			38404: outdata = 32'd27132;
			38405: outdata = 32'd27131;
			38406: outdata = 32'd27130;
			38407: outdata = 32'd27129;
			38408: outdata = 32'd27128;
			38409: outdata = 32'd27127;
			38410: outdata = 32'd27126;
			38411: outdata = 32'd27125;
			38412: outdata = 32'd27124;
			38413: outdata = 32'd27123;
			38414: outdata = 32'd27122;
			38415: outdata = 32'd27121;
			38416: outdata = 32'd27120;
			38417: outdata = 32'd27119;
			38418: outdata = 32'd27118;
			38419: outdata = 32'd27117;
			38420: outdata = 32'd27116;
			38421: outdata = 32'd27115;
			38422: outdata = 32'd27114;
			38423: outdata = 32'd27113;
			38424: outdata = 32'd27112;
			38425: outdata = 32'd27111;
			38426: outdata = 32'd27110;
			38427: outdata = 32'd27109;
			38428: outdata = 32'd27108;
			38429: outdata = 32'd27107;
			38430: outdata = 32'd27106;
			38431: outdata = 32'd27105;
			38432: outdata = 32'd27104;
			38433: outdata = 32'd27103;
			38434: outdata = 32'd27102;
			38435: outdata = 32'd27101;
			38436: outdata = 32'd27100;
			38437: outdata = 32'd27099;
			38438: outdata = 32'd27098;
			38439: outdata = 32'd27097;
			38440: outdata = 32'd27096;
			38441: outdata = 32'd27095;
			38442: outdata = 32'd27094;
			38443: outdata = 32'd27093;
			38444: outdata = 32'd27092;
			38445: outdata = 32'd27091;
			38446: outdata = 32'd27090;
			38447: outdata = 32'd27089;
			38448: outdata = 32'd27088;
			38449: outdata = 32'd27087;
			38450: outdata = 32'd27086;
			38451: outdata = 32'd27085;
			38452: outdata = 32'd27084;
			38453: outdata = 32'd27083;
			38454: outdata = 32'd27082;
			38455: outdata = 32'd27081;
			38456: outdata = 32'd27080;
			38457: outdata = 32'd27079;
			38458: outdata = 32'd27078;
			38459: outdata = 32'd27077;
			38460: outdata = 32'd27076;
			38461: outdata = 32'd27075;
			38462: outdata = 32'd27074;
			38463: outdata = 32'd27073;
			38464: outdata = 32'd27072;
			38465: outdata = 32'd27071;
			38466: outdata = 32'd27070;
			38467: outdata = 32'd27069;
			38468: outdata = 32'd27068;
			38469: outdata = 32'd27067;
			38470: outdata = 32'd27066;
			38471: outdata = 32'd27065;
			38472: outdata = 32'd27064;
			38473: outdata = 32'd27063;
			38474: outdata = 32'd27062;
			38475: outdata = 32'd27061;
			38476: outdata = 32'd27060;
			38477: outdata = 32'd27059;
			38478: outdata = 32'd27058;
			38479: outdata = 32'd27057;
			38480: outdata = 32'd27056;
			38481: outdata = 32'd27055;
			38482: outdata = 32'd27054;
			38483: outdata = 32'd27053;
			38484: outdata = 32'd27052;
			38485: outdata = 32'd27051;
			38486: outdata = 32'd27050;
			38487: outdata = 32'd27049;
			38488: outdata = 32'd27048;
			38489: outdata = 32'd27047;
			38490: outdata = 32'd27046;
			38491: outdata = 32'd27045;
			38492: outdata = 32'd27044;
			38493: outdata = 32'd27043;
			38494: outdata = 32'd27042;
			38495: outdata = 32'd27041;
			38496: outdata = 32'd27040;
			38497: outdata = 32'd27039;
			38498: outdata = 32'd27038;
			38499: outdata = 32'd27037;
			38500: outdata = 32'd27036;
			38501: outdata = 32'd27035;
			38502: outdata = 32'd27034;
			38503: outdata = 32'd27033;
			38504: outdata = 32'd27032;
			38505: outdata = 32'd27031;
			38506: outdata = 32'd27030;
			38507: outdata = 32'd27029;
			38508: outdata = 32'd27028;
			38509: outdata = 32'd27027;
			38510: outdata = 32'd27026;
			38511: outdata = 32'd27025;
			38512: outdata = 32'd27024;
			38513: outdata = 32'd27023;
			38514: outdata = 32'd27022;
			38515: outdata = 32'd27021;
			38516: outdata = 32'd27020;
			38517: outdata = 32'd27019;
			38518: outdata = 32'd27018;
			38519: outdata = 32'd27017;
			38520: outdata = 32'd27016;
			38521: outdata = 32'd27015;
			38522: outdata = 32'd27014;
			38523: outdata = 32'd27013;
			38524: outdata = 32'd27012;
			38525: outdata = 32'd27011;
			38526: outdata = 32'd27010;
			38527: outdata = 32'd27009;
			38528: outdata = 32'd27008;
			38529: outdata = 32'd27007;
			38530: outdata = 32'd27006;
			38531: outdata = 32'd27005;
			38532: outdata = 32'd27004;
			38533: outdata = 32'd27003;
			38534: outdata = 32'd27002;
			38535: outdata = 32'd27001;
			38536: outdata = 32'd27000;
			38537: outdata = 32'd26999;
			38538: outdata = 32'd26998;
			38539: outdata = 32'd26997;
			38540: outdata = 32'd26996;
			38541: outdata = 32'd26995;
			38542: outdata = 32'd26994;
			38543: outdata = 32'd26993;
			38544: outdata = 32'd26992;
			38545: outdata = 32'd26991;
			38546: outdata = 32'd26990;
			38547: outdata = 32'd26989;
			38548: outdata = 32'd26988;
			38549: outdata = 32'd26987;
			38550: outdata = 32'd26986;
			38551: outdata = 32'd26985;
			38552: outdata = 32'd26984;
			38553: outdata = 32'd26983;
			38554: outdata = 32'd26982;
			38555: outdata = 32'd26981;
			38556: outdata = 32'd26980;
			38557: outdata = 32'd26979;
			38558: outdata = 32'd26978;
			38559: outdata = 32'd26977;
			38560: outdata = 32'd26976;
			38561: outdata = 32'd26975;
			38562: outdata = 32'd26974;
			38563: outdata = 32'd26973;
			38564: outdata = 32'd26972;
			38565: outdata = 32'd26971;
			38566: outdata = 32'd26970;
			38567: outdata = 32'd26969;
			38568: outdata = 32'd26968;
			38569: outdata = 32'd26967;
			38570: outdata = 32'd26966;
			38571: outdata = 32'd26965;
			38572: outdata = 32'd26964;
			38573: outdata = 32'd26963;
			38574: outdata = 32'd26962;
			38575: outdata = 32'd26961;
			38576: outdata = 32'd26960;
			38577: outdata = 32'd26959;
			38578: outdata = 32'd26958;
			38579: outdata = 32'd26957;
			38580: outdata = 32'd26956;
			38581: outdata = 32'd26955;
			38582: outdata = 32'd26954;
			38583: outdata = 32'd26953;
			38584: outdata = 32'd26952;
			38585: outdata = 32'd26951;
			38586: outdata = 32'd26950;
			38587: outdata = 32'd26949;
			38588: outdata = 32'd26948;
			38589: outdata = 32'd26947;
			38590: outdata = 32'd26946;
			38591: outdata = 32'd26945;
			38592: outdata = 32'd26944;
			38593: outdata = 32'd26943;
			38594: outdata = 32'd26942;
			38595: outdata = 32'd26941;
			38596: outdata = 32'd26940;
			38597: outdata = 32'd26939;
			38598: outdata = 32'd26938;
			38599: outdata = 32'd26937;
			38600: outdata = 32'd26936;
			38601: outdata = 32'd26935;
			38602: outdata = 32'd26934;
			38603: outdata = 32'd26933;
			38604: outdata = 32'd26932;
			38605: outdata = 32'd26931;
			38606: outdata = 32'd26930;
			38607: outdata = 32'd26929;
			38608: outdata = 32'd26928;
			38609: outdata = 32'd26927;
			38610: outdata = 32'd26926;
			38611: outdata = 32'd26925;
			38612: outdata = 32'd26924;
			38613: outdata = 32'd26923;
			38614: outdata = 32'd26922;
			38615: outdata = 32'd26921;
			38616: outdata = 32'd26920;
			38617: outdata = 32'd26919;
			38618: outdata = 32'd26918;
			38619: outdata = 32'd26917;
			38620: outdata = 32'd26916;
			38621: outdata = 32'd26915;
			38622: outdata = 32'd26914;
			38623: outdata = 32'd26913;
			38624: outdata = 32'd26912;
			38625: outdata = 32'd26911;
			38626: outdata = 32'd26910;
			38627: outdata = 32'd26909;
			38628: outdata = 32'd26908;
			38629: outdata = 32'd26907;
			38630: outdata = 32'd26906;
			38631: outdata = 32'd26905;
			38632: outdata = 32'd26904;
			38633: outdata = 32'd26903;
			38634: outdata = 32'd26902;
			38635: outdata = 32'd26901;
			38636: outdata = 32'd26900;
			38637: outdata = 32'd26899;
			38638: outdata = 32'd26898;
			38639: outdata = 32'd26897;
			38640: outdata = 32'd26896;
			38641: outdata = 32'd26895;
			38642: outdata = 32'd26894;
			38643: outdata = 32'd26893;
			38644: outdata = 32'd26892;
			38645: outdata = 32'd26891;
			38646: outdata = 32'd26890;
			38647: outdata = 32'd26889;
			38648: outdata = 32'd26888;
			38649: outdata = 32'd26887;
			38650: outdata = 32'd26886;
			38651: outdata = 32'd26885;
			38652: outdata = 32'd26884;
			38653: outdata = 32'd26883;
			38654: outdata = 32'd26882;
			38655: outdata = 32'd26881;
			38656: outdata = 32'd26880;
			38657: outdata = 32'd26879;
			38658: outdata = 32'd26878;
			38659: outdata = 32'd26877;
			38660: outdata = 32'd26876;
			38661: outdata = 32'd26875;
			38662: outdata = 32'd26874;
			38663: outdata = 32'd26873;
			38664: outdata = 32'd26872;
			38665: outdata = 32'd26871;
			38666: outdata = 32'd26870;
			38667: outdata = 32'd26869;
			38668: outdata = 32'd26868;
			38669: outdata = 32'd26867;
			38670: outdata = 32'd26866;
			38671: outdata = 32'd26865;
			38672: outdata = 32'd26864;
			38673: outdata = 32'd26863;
			38674: outdata = 32'd26862;
			38675: outdata = 32'd26861;
			38676: outdata = 32'd26860;
			38677: outdata = 32'd26859;
			38678: outdata = 32'd26858;
			38679: outdata = 32'd26857;
			38680: outdata = 32'd26856;
			38681: outdata = 32'd26855;
			38682: outdata = 32'd26854;
			38683: outdata = 32'd26853;
			38684: outdata = 32'd26852;
			38685: outdata = 32'd26851;
			38686: outdata = 32'd26850;
			38687: outdata = 32'd26849;
			38688: outdata = 32'd26848;
			38689: outdata = 32'd26847;
			38690: outdata = 32'd26846;
			38691: outdata = 32'd26845;
			38692: outdata = 32'd26844;
			38693: outdata = 32'd26843;
			38694: outdata = 32'd26842;
			38695: outdata = 32'd26841;
			38696: outdata = 32'd26840;
			38697: outdata = 32'd26839;
			38698: outdata = 32'd26838;
			38699: outdata = 32'd26837;
			38700: outdata = 32'd26836;
			38701: outdata = 32'd26835;
			38702: outdata = 32'd26834;
			38703: outdata = 32'd26833;
			38704: outdata = 32'd26832;
			38705: outdata = 32'd26831;
			38706: outdata = 32'd26830;
			38707: outdata = 32'd26829;
			38708: outdata = 32'd26828;
			38709: outdata = 32'd26827;
			38710: outdata = 32'd26826;
			38711: outdata = 32'd26825;
			38712: outdata = 32'd26824;
			38713: outdata = 32'd26823;
			38714: outdata = 32'd26822;
			38715: outdata = 32'd26821;
			38716: outdata = 32'd26820;
			38717: outdata = 32'd26819;
			38718: outdata = 32'd26818;
			38719: outdata = 32'd26817;
			38720: outdata = 32'd26816;
			38721: outdata = 32'd26815;
			38722: outdata = 32'd26814;
			38723: outdata = 32'd26813;
			38724: outdata = 32'd26812;
			38725: outdata = 32'd26811;
			38726: outdata = 32'd26810;
			38727: outdata = 32'd26809;
			38728: outdata = 32'd26808;
			38729: outdata = 32'd26807;
			38730: outdata = 32'd26806;
			38731: outdata = 32'd26805;
			38732: outdata = 32'd26804;
			38733: outdata = 32'd26803;
			38734: outdata = 32'd26802;
			38735: outdata = 32'd26801;
			38736: outdata = 32'd26800;
			38737: outdata = 32'd26799;
			38738: outdata = 32'd26798;
			38739: outdata = 32'd26797;
			38740: outdata = 32'd26796;
			38741: outdata = 32'd26795;
			38742: outdata = 32'd26794;
			38743: outdata = 32'd26793;
			38744: outdata = 32'd26792;
			38745: outdata = 32'd26791;
			38746: outdata = 32'd26790;
			38747: outdata = 32'd26789;
			38748: outdata = 32'd26788;
			38749: outdata = 32'd26787;
			38750: outdata = 32'd26786;
			38751: outdata = 32'd26785;
			38752: outdata = 32'd26784;
			38753: outdata = 32'd26783;
			38754: outdata = 32'd26782;
			38755: outdata = 32'd26781;
			38756: outdata = 32'd26780;
			38757: outdata = 32'd26779;
			38758: outdata = 32'd26778;
			38759: outdata = 32'd26777;
			38760: outdata = 32'd26776;
			38761: outdata = 32'd26775;
			38762: outdata = 32'd26774;
			38763: outdata = 32'd26773;
			38764: outdata = 32'd26772;
			38765: outdata = 32'd26771;
			38766: outdata = 32'd26770;
			38767: outdata = 32'd26769;
			38768: outdata = 32'd26768;
			38769: outdata = 32'd26767;
			38770: outdata = 32'd26766;
			38771: outdata = 32'd26765;
			38772: outdata = 32'd26764;
			38773: outdata = 32'd26763;
			38774: outdata = 32'd26762;
			38775: outdata = 32'd26761;
			38776: outdata = 32'd26760;
			38777: outdata = 32'd26759;
			38778: outdata = 32'd26758;
			38779: outdata = 32'd26757;
			38780: outdata = 32'd26756;
			38781: outdata = 32'd26755;
			38782: outdata = 32'd26754;
			38783: outdata = 32'd26753;
			38784: outdata = 32'd26752;
			38785: outdata = 32'd26751;
			38786: outdata = 32'd26750;
			38787: outdata = 32'd26749;
			38788: outdata = 32'd26748;
			38789: outdata = 32'd26747;
			38790: outdata = 32'd26746;
			38791: outdata = 32'd26745;
			38792: outdata = 32'd26744;
			38793: outdata = 32'd26743;
			38794: outdata = 32'd26742;
			38795: outdata = 32'd26741;
			38796: outdata = 32'd26740;
			38797: outdata = 32'd26739;
			38798: outdata = 32'd26738;
			38799: outdata = 32'd26737;
			38800: outdata = 32'd26736;
			38801: outdata = 32'd26735;
			38802: outdata = 32'd26734;
			38803: outdata = 32'd26733;
			38804: outdata = 32'd26732;
			38805: outdata = 32'd26731;
			38806: outdata = 32'd26730;
			38807: outdata = 32'd26729;
			38808: outdata = 32'd26728;
			38809: outdata = 32'd26727;
			38810: outdata = 32'd26726;
			38811: outdata = 32'd26725;
			38812: outdata = 32'd26724;
			38813: outdata = 32'd26723;
			38814: outdata = 32'd26722;
			38815: outdata = 32'd26721;
			38816: outdata = 32'd26720;
			38817: outdata = 32'd26719;
			38818: outdata = 32'd26718;
			38819: outdata = 32'd26717;
			38820: outdata = 32'd26716;
			38821: outdata = 32'd26715;
			38822: outdata = 32'd26714;
			38823: outdata = 32'd26713;
			38824: outdata = 32'd26712;
			38825: outdata = 32'd26711;
			38826: outdata = 32'd26710;
			38827: outdata = 32'd26709;
			38828: outdata = 32'd26708;
			38829: outdata = 32'd26707;
			38830: outdata = 32'd26706;
			38831: outdata = 32'd26705;
			38832: outdata = 32'd26704;
			38833: outdata = 32'd26703;
			38834: outdata = 32'd26702;
			38835: outdata = 32'd26701;
			38836: outdata = 32'd26700;
			38837: outdata = 32'd26699;
			38838: outdata = 32'd26698;
			38839: outdata = 32'd26697;
			38840: outdata = 32'd26696;
			38841: outdata = 32'd26695;
			38842: outdata = 32'd26694;
			38843: outdata = 32'd26693;
			38844: outdata = 32'd26692;
			38845: outdata = 32'd26691;
			38846: outdata = 32'd26690;
			38847: outdata = 32'd26689;
			38848: outdata = 32'd26688;
			38849: outdata = 32'd26687;
			38850: outdata = 32'd26686;
			38851: outdata = 32'd26685;
			38852: outdata = 32'd26684;
			38853: outdata = 32'd26683;
			38854: outdata = 32'd26682;
			38855: outdata = 32'd26681;
			38856: outdata = 32'd26680;
			38857: outdata = 32'd26679;
			38858: outdata = 32'd26678;
			38859: outdata = 32'd26677;
			38860: outdata = 32'd26676;
			38861: outdata = 32'd26675;
			38862: outdata = 32'd26674;
			38863: outdata = 32'd26673;
			38864: outdata = 32'd26672;
			38865: outdata = 32'd26671;
			38866: outdata = 32'd26670;
			38867: outdata = 32'd26669;
			38868: outdata = 32'd26668;
			38869: outdata = 32'd26667;
			38870: outdata = 32'd26666;
			38871: outdata = 32'd26665;
			38872: outdata = 32'd26664;
			38873: outdata = 32'd26663;
			38874: outdata = 32'd26662;
			38875: outdata = 32'd26661;
			38876: outdata = 32'd26660;
			38877: outdata = 32'd26659;
			38878: outdata = 32'd26658;
			38879: outdata = 32'd26657;
			38880: outdata = 32'd26656;
			38881: outdata = 32'd26655;
			38882: outdata = 32'd26654;
			38883: outdata = 32'd26653;
			38884: outdata = 32'd26652;
			38885: outdata = 32'd26651;
			38886: outdata = 32'd26650;
			38887: outdata = 32'd26649;
			38888: outdata = 32'd26648;
			38889: outdata = 32'd26647;
			38890: outdata = 32'd26646;
			38891: outdata = 32'd26645;
			38892: outdata = 32'd26644;
			38893: outdata = 32'd26643;
			38894: outdata = 32'd26642;
			38895: outdata = 32'd26641;
			38896: outdata = 32'd26640;
			38897: outdata = 32'd26639;
			38898: outdata = 32'd26638;
			38899: outdata = 32'd26637;
			38900: outdata = 32'd26636;
			38901: outdata = 32'd26635;
			38902: outdata = 32'd26634;
			38903: outdata = 32'd26633;
			38904: outdata = 32'd26632;
			38905: outdata = 32'd26631;
			38906: outdata = 32'd26630;
			38907: outdata = 32'd26629;
			38908: outdata = 32'd26628;
			38909: outdata = 32'd26627;
			38910: outdata = 32'd26626;
			38911: outdata = 32'd26625;
			38912: outdata = 32'd26624;
			38913: outdata = 32'd26623;
			38914: outdata = 32'd26622;
			38915: outdata = 32'd26621;
			38916: outdata = 32'd26620;
			38917: outdata = 32'd26619;
			38918: outdata = 32'd26618;
			38919: outdata = 32'd26617;
			38920: outdata = 32'd26616;
			38921: outdata = 32'd26615;
			38922: outdata = 32'd26614;
			38923: outdata = 32'd26613;
			38924: outdata = 32'd26612;
			38925: outdata = 32'd26611;
			38926: outdata = 32'd26610;
			38927: outdata = 32'd26609;
			38928: outdata = 32'd26608;
			38929: outdata = 32'd26607;
			38930: outdata = 32'd26606;
			38931: outdata = 32'd26605;
			38932: outdata = 32'd26604;
			38933: outdata = 32'd26603;
			38934: outdata = 32'd26602;
			38935: outdata = 32'd26601;
			38936: outdata = 32'd26600;
			38937: outdata = 32'd26599;
			38938: outdata = 32'd26598;
			38939: outdata = 32'd26597;
			38940: outdata = 32'd26596;
			38941: outdata = 32'd26595;
			38942: outdata = 32'd26594;
			38943: outdata = 32'd26593;
			38944: outdata = 32'd26592;
			38945: outdata = 32'd26591;
			38946: outdata = 32'd26590;
			38947: outdata = 32'd26589;
			38948: outdata = 32'd26588;
			38949: outdata = 32'd26587;
			38950: outdata = 32'd26586;
			38951: outdata = 32'd26585;
			38952: outdata = 32'd26584;
			38953: outdata = 32'd26583;
			38954: outdata = 32'd26582;
			38955: outdata = 32'd26581;
			38956: outdata = 32'd26580;
			38957: outdata = 32'd26579;
			38958: outdata = 32'd26578;
			38959: outdata = 32'd26577;
			38960: outdata = 32'd26576;
			38961: outdata = 32'd26575;
			38962: outdata = 32'd26574;
			38963: outdata = 32'd26573;
			38964: outdata = 32'd26572;
			38965: outdata = 32'd26571;
			38966: outdata = 32'd26570;
			38967: outdata = 32'd26569;
			38968: outdata = 32'd26568;
			38969: outdata = 32'd26567;
			38970: outdata = 32'd26566;
			38971: outdata = 32'd26565;
			38972: outdata = 32'd26564;
			38973: outdata = 32'd26563;
			38974: outdata = 32'd26562;
			38975: outdata = 32'd26561;
			38976: outdata = 32'd26560;
			38977: outdata = 32'd26559;
			38978: outdata = 32'd26558;
			38979: outdata = 32'd26557;
			38980: outdata = 32'd26556;
			38981: outdata = 32'd26555;
			38982: outdata = 32'd26554;
			38983: outdata = 32'd26553;
			38984: outdata = 32'd26552;
			38985: outdata = 32'd26551;
			38986: outdata = 32'd26550;
			38987: outdata = 32'd26549;
			38988: outdata = 32'd26548;
			38989: outdata = 32'd26547;
			38990: outdata = 32'd26546;
			38991: outdata = 32'd26545;
			38992: outdata = 32'd26544;
			38993: outdata = 32'd26543;
			38994: outdata = 32'd26542;
			38995: outdata = 32'd26541;
			38996: outdata = 32'd26540;
			38997: outdata = 32'd26539;
			38998: outdata = 32'd26538;
			38999: outdata = 32'd26537;
			39000: outdata = 32'd26536;
			39001: outdata = 32'd26535;
			39002: outdata = 32'd26534;
			39003: outdata = 32'd26533;
			39004: outdata = 32'd26532;
			39005: outdata = 32'd26531;
			39006: outdata = 32'd26530;
			39007: outdata = 32'd26529;
			39008: outdata = 32'd26528;
			39009: outdata = 32'd26527;
			39010: outdata = 32'd26526;
			39011: outdata = 32'd26525;
			39012: outdata = 32'd26524;
			39013: outdata = 32'd26523;
			39014: outdata = 32'd26522;
			39015: outdata = 32'd26521;
			39016: outdata = 32'd26520;
			39017: outdata = 32'd26519;
			39018: outdata = 32'd26518;
			39019: outdata = 32'd26517;
			39020: outdata = 32'd26516;
			39021: outdata = 32'd26515;
			39022: outdata = 32'd26514;
			39023: outdata = 32'd26513;
			39024: outdata = 32'd26512;
			39025: outdata = 32'd26511;
			39026: outdata = 32'd26510;
			39027: outdata = 32'd26509;
			39028: outdata = 32'd26508;
			39029: outdata = 32'd26507;
			39030: outdata = 32'd26506;
			39031: outdata = 32'd26505;
			39032: outdata = 32'd26504;
			39033: outdata = 32'd26503;
			39034: outdata = 32'd26502;
			39035: outdata = 32'd26501;
			39036: outdata = 32'd26500;
			39037: outdata = 32'd26499;
			39038: outdata = 32'd26498;
			39039: outdata = 32'd26497;
			39040: outdata = 32'd26496;
			39041: outdata = 32'd26495;
			39042: outdata = 32'd26494;
			39043: outdata = 32'd26493;
			39044: outdata = 32'd26492;
			39045: outdata = 32'd26491;
			39046: outdata = 32'd26490;
			39047: outdata = 32'd26489;
			39048: outdata = 32'd26488;
			39049: outdata = 32'd26487;
			39050: outdata = 32'd26486;
			39051: outdata = 32'd26485;
			39052: outdata = 32'd26484;
			39053: outdata = 32'd26483;
			39054: outdata = 32'd26482;
			39055: outdata = 32'd26481;
			39056: outdata = 32'd26480;
			39057: outdata = 32'd26479;
			39058: outdata = 32'd26478;
			39059: outdata = 32'd26477;
			39060: outdata = 32'd26476;
			39061: outdata = 32'd26475;
			39062: outdata = 32'd26474;
			39063: outdata = 32'd26473;
			39064: outdata = 32'd26472;
			39065: outdata = 32'd26471;
			39066: outdata = 32'd26470;
			39067: outdata = 32'd26469;
			39068: outdata = 32'd26468;
			39069: outdata = 32'd26467;
			39070: outdata = 32'd26466;
			39071: outdata = 32'd26465;
			39072: outdata = 32'd26464;
			39073: outdata = 32'd26463;
			39074: outdata = 32'd26462;
			39075: outdata = 32'd26461;
			39076: outdata = 32'd26460;
			39077: outdata = 32'd26459;
			39078: outdata = 32'd26458;
			39079: outdata = 32'd26457;
			39080: outdata = 32'd26456;
			39081: outdata = 32'd26455;
			39082: outdata = 32'd26454;
			39083: outdata = 32'd26453;
			39084: outdata = 32'd26452;
			39085: outdata = 32'd26451;
			39086: outdata = 32'd26450;
			39087: outdata = 32'd26449;
			39088: outdata = 32'd26448;
			39089: outdata = 32'd26447;
			39090: outdata = 32'd26446;
			39091: outdata = 32'd26445;
			39092: outdata = 32'd26444;
			39093: outdata = 32'd26443;
			39094: outdata = 32'd26442;
			39095: outdata = 32'd26441;
			39096: outdata = 32'd26440;
			39097: outdata = 32'd26439;
			39098: outdata = 32'd26438;
			39099: outdata = 32'd26437;
			39100: outdata = 32'd26436;
			39101: outdata = 32'd26435;
			39102: outdata = 32'd26434;
			39103: outdata = 32'd26433;
			39104: outdata = 32'd26432;
			39105: outdata = 32'd26431;
			39106: outdata = 32'd26430;
			39107: outdata = 32'd26429;
			39108: outdata = 32'd26428;
			39109: outdata = 32'd26427;
			39110: outdata = 32'd26426;
			39111: outdata = 32'd26425;
			39112: outdata = 32'd26424;
			39113: outdata = 32'd26423;
			39114: outdata = 32'd26422;
			39115: outdata = 32'd26421;
			39116: outdata = 32'd26420;
			39117: outdata = 32'd26419;
			39118: outdata = 32'd26418;
			39119: outdata = 32'd26417;
			39120: outdata = 32'd26416;
			39121: outdata = 32'd26415;
			39122: outdata = 32'd26414;
			39123: outdata = 32'd26413;
			39124: outdata = 32'd26412;
			39125: outdata = 32'd26411;
			39126: outdata = 32'd26410;
			39127: outdata = 32'd26409;
			39128: outdata = 32'd26408;
			39129: outdata = 32'd26407;
			39130: outdata = 32'd26406;
			39131: outdata = 32'd26405;
			39132: outdata = 32'd26404;
			39133: outdata = 32'd26403;
			39134: outdata = 32'd26402;
			39135: outdata = 32'd26401;
			39136: outdata = 32'd26400;
			39137: outdata = 32'd26399;
			39138: outdata = 32'd26398;
			39139: outdata = 32'd26397;
			39140: outdata = 32'd26396;
			39141: outdata = 32'd26395;
			39142: outdata = 32'd26394;
			39143: outdata = 32'd26393;
			39144: outdata = 32'd26392;
			39145: outdata = 32'd26391;
			39146: outdata = 32'd26390;
			39147: outdata = 32'd26389;
			39148: outdata = 32'd26388;
			39149: outdata = 32'd26387;
			39150: outdata = 32'd26386;
			39151: outdata = 32'd26385;
			39152: outdata = 32'd26384;
			39153: outdata = 32'd26383;
			39154: outdata = 32'd26382;
			39155: outdata = 32'd26381;
			39156: outdata = 32'd26380;
			39157: outdata = 32'd26379;
			39158: outdata = 32'd26378;
			39159: outdata = 32'd26377;
			39160: outdata = 32'd26376;
			39161: outdata = 32'd26375;
			39162: outdata = 32'd26374;
			39163: outdata = 32'd26373;
			39164: outdata = 32'd26372;
			39165: outdata = 32'd26371;
			39166: outdata = 32'd26370;
			39167: outdata = 32'd26369;
			39168: outdata = 32'd26368;
			39169: outdata = 32'd26367;
			39170: outdata = 32'd26366;
			39171: outdata = 32'd26365;
			39172: outdata = 32'd26364;
			39173: outdata = 32'd26363;
			39174: outdata = 32'd26362;
			39175: outdata = 32'd26361;
			39176: outdata = 32'd26360;
			39177: outdata = 32'd26359;
			39178: outdata = 32'd26358;
			39179: outdata = 32'd26357;
			39180: outdata = 32'd26356;
			39181: outdata = 32'd26355;
			39182: outdata = 32'd26354;
			39183: outdata = 32'd26353;
			39184: outdata = 32'd26352;
			39185: outdata = 32'd26351;
			39186: outdata = 32'd26350;
			39187: outdata = 32'd26349;
			39188: outdata = 32'd26348;
			39189: outdata = 32'd26347;
			39190: outdata = 32'd26346;
			39191: outdata = 32'd26345;
			39192: outdata = 32'd26344;
			39193: outdata = 32'd26343;
			39194: outdata = 32'd26342;
			39195: outdata = 32'd26341;
			39196: outdata = 32'd26340;
			39197: outdata = 32'd26339;
			39198: outdata = 32'd26338;
			39199: outdata = 32'd26337;
			39200: outdata = 32'd26336;
			39201: outdata = 32'd26335;
			39202: outdata = 32'd26334;
			39203: outdata = 32'd26333;
			39204: outdata = 32'd26332;
			39205: outdata = 32'd26331;
			39206: outdata = 32'd26330;
			39207: outdata = 32'd26329;
			39208: outdata = 32'd26328;
			39209: outdata = 32'd26327;
			39210: outdata = 32'd26326;
			39211: outdata = 32'd26325;
			39212: outdata = 32'd26324;
			39213: outdata = 32'd26323;
			39214: outdata = 32'd26322;
			39215: outdata = 32'd26321;
			39216: outdata = 32'd26320;
			39217: outdata = 32'd26319;
			39218: outdata = 32'd26318;
			39219: outdata = 32'd26317;
			39220: outdata = 32'd26316;
			39221: outdata = 32'd26315;
			39222: outdata = 32'd26314;
			39223: outdata = 32'd26313;
			39224: outdata = 32'd26312;
			39225: outdata = 32'd26311;
			39226: outdata = 32'd26310;
			39227: outdata = 32'd26309;
			39228: outdata = 32'd26308;
			39229: outdata = 32'd26307;
			39230: outdata = 32'd26306;
			39231: outdata = 32'd26305;
			39232: outdata = 32'd26304;
			39233: outdata = 32'd26303;
			39234: outdata = 32'd26302;
			39235: outdata = 32'd26301;
			39236: outdata = 32'd26300;
			39237: outdata = 32'd26299;
			39238: outdata = 32'd26298;
			39239: outdata = 32'd26297;
			39240: outdata = 32'd26296;
			39241: outdata = 32'd26295;
			39242: outdata = 32'd26294;
			39243: outdata = 32'd26293;
			39244: outdata = 32'd26292;
			39245: outdata = 32'd26291;
			39246: outdata = 32'd26290;
			39247: outdata = 32'd26289;
			39248: outdata = 32'd26288;
			39249: outdata = 32'd26287;
			39250: outdata = 32'd26286;
			39251: outdata = 32'd26285;
			39252: outdata = 32'd26284;
			39253: outdata = 32'd26283;
			39254: outdata = 32'd26282;
			39255: outdata = 32'd26281;
			39256: outdata = 32'd26280;
			39257: outdata = 32'd26279;
			39258: outdata = 32'd26278;
			39259: outdata = 32'd26277;
			39260: outdata = 32'd26276;
			39261: outdata = 32'd26275;
			39262: outdata = 32'd26274;
			39263: outdata = 32'd26273;
			39264: outdata = 32'd26272;
			39265: outdata = 32'd26271;
			39266: outdata = 32'd26270;
			39267: outdata = 32'd26269;
			39268: outdata = 32'd26268;
			39269: outdata = 32'd26267;
			39270: outdata = 32'd26266;
			39271: outdata = 32'd26265;
			39272: outdata = 32'd26264;
			39273: outdata = 32'd26263;
			39274: outdata = 32'd26262;
			39275: outdata = 32'd26261;
			39276: outdata = 32'd26260;
			39277: outdata = 32'd26259;
			39278: outdata = 32'd26258;
			39279: outdata = 32'd26257;
			39280: outdata = 32'd26256;
			39281: outdata = 32'd26255;
			39282: outdata = 32'd26254;
			39283: outdata = 32'd26253;
			39284: outdata = 32'd26252;
			39285: outdata = 32'd26251;
			39286: outdata = 32'd26250;
			39287: outdata = 32'd26249;
			39288: outdata = 32'd26248;
			39289: outdata = 32'd26247;
			39290: outdata = 32'd26246;
			39291: outdata = 32'd26245;
			39292: outdata = 32'd26244;
			39293: outdata = 32'd26243;
			39294: outdata = 32'd26242;
			39295: outdata = 32'd26241;
			39296: outdata = 32'd26240;
			39297: outdata = 32'd26239;
			39298: outdata = 32'd26238;
			39299: outdata = 32'd26237;
			39300: outdata = 32'd26236;
			39301: outdata = 32'd26235;
			39302: outdata = 32'd26234;
			39303: outdata = 32'd26233;
			39304: outdata = 32'd26232;
			39305: outdata = 32'd26231;
			39306: outdata = 32'd26230;
			39307: outdata = 32'd26229;
			39308: outdata = 32'd26228;
			39309: outdata = 32'd26227;
			39310: outdata = 32'd26226;
			39311: outdata = 32'd26225;
			39312: outdata = 32'd26224;
			39313: outdata = 32'd26223;
			39314: outdata = 32'd26222;
			39315: outdata = 32'd26221;
			39316: outdata = 32'd26220;
			39317: outdata = 32'd26219;
			39318: outdata = 32'd26218;
			39319: outdata = 32'd26217;
			39320: outdata = 32'd26216;
			39321: outdata = 32'd26215;
			39322: outdata = 32'd26214;
			39323: outdata = 32'd26213;
			39324: outdata = 32'd26212;
			39325: outdata = 32'd26211;
			39326: outdata = 32'd26210;
			39327: outdata = 32'd26209;
			39328: outdata = 32'd26208;
			39329: outdata = 32'd26207;
			39330: outdata = 32'd26206;
			39331: outdata = 32'd26205;
			39332: outdata = 32'd26204;
			39333: outdata = 32'd26203;
			39334: outdata = 32'd26202;
			39335: outdata = 32'd26201;
			39336: outdata = 32'd26200;
			39337: outdata = 32'd26199;
			39338: outdata = 32'd26198;
			39339: outdata = 32'd26197;
			39340: outdata = 32'd26196;
			39341: outdata = 32'd26195;
			39342: outdata = 32'd26194;
			39343: outdata = 32'd26193;
			39344: outdata = 32'd26192;
			39345: outdata = 32'd26191;
			39346: outdata = 32'd26190;
			39347: outdata = 32'd26189;
			39348: outdata = 32'd26188;
			39349: outdata = 32'd26187;
			39350: outdata = 32'd26186;
			39351: outdata = 32'd26185;
			39352: outdata = 32'd26184;
			39353: outdata = 32'd26183;
			39354: outdata = 32'd26182;
			39355: outdata = 32'd26181;
			39356: outdata = 32'd26180;
			39357: outdata = 32'd26179;
			39358: outdata = 32'd26178;
			39359: outdata = 32'd26177;
			39360: outdata = 32'd26176;
			39361: outdata = 32'd26175;
			39362: outdata = 32'd26174;
			39363: outdata = 32'd26173;
			39364: outdata = 32'd26172;
			39365: outdata = 32'd26171;
			39366: outdata = 32'd26170;
			39367: outdata = 32'd26169;
			39368: outdata = 32'd26168;
			39369: outdata = 32'd26167;
			39370: outdata = 32'd26166;
			39371: outdata = 32'd26165;
			39372: outdata = 32'd26164;
			39373: outdata = 32'd26163;
			39374: outdata = 32'd26162;
			39375: outdata = 32'd26161;
			39376: outdata = 32'd26160;
			39377: outdata = 32'd26159;
			39378: outdata = 32'd26158;
			39379: outdata = 32'd26157;
			39380: outdata = 32'd26156;
			39381: outdata = 32'd26155;
			39382: outdata = 32'd26154;
			39383: outdata = 32'd26153;
			39384: outdata = 32'd26152;
			39385: outdata = 32'd26151;
			39386: outdata = 32'd26150;
			39387: outdata = 32'd26149;
			39388: outdata = 32'd26148;
			39389: outdata = 32'd26147;
			39390: outdata = 32'd26146;
			39391: outdata = 32'd26145;
			39392: outdata = 32'd26144;
			39393: outdata = 32'd26143;
			39394: outdata = 32'd26142;
			39395: outdata = 32'd26141;
			39396: outdata = 32'd26140;
			39397: outdata = 32'd26139;
			39398: outdata = 32'd26138;
			39399: outdata = 32'd26137;
			39400: outdata = 32'd26136;
			39401: outdata = 32'd26135;
			39402: outdata = 32'd26134;
			39403: outdata = 32'd26133;
			39404: outdata = 32'd26132;
			39405: outdata = 32'd26131;
			39406: outdata = 32'd26130;
			39407: outdata = 32'd26129;
			39408: outdata = 32'd26128;
			39409: outdata = 32'd26127;
			39410: outdata = 32'd26126;
			39411: outdata = 32'd26125;
			39412: outdata = 32'd26124;
			39413: outdata = 32'd26123;
			39414: outdata = 32'd26122;
			39415: outdata = 32'd26121;
			39416: outdata = 32'd26120;
			39417: outdata = 32'd26119;
			39418: outdata = 32'd26118;
			39419: outdata = 32'd26117;
			39420: outdata = 32'd26116;
			39421: outdata = 32'd26115;
			39422: outdata = 32'd26114;
			39423: outdata = 32'd26113;
			39424: outdata = 32'd26112;
			39425: outdata = 32'd26111;
			39426: outdata = 32'd26110;
			39427: outdata = 32'd26109;
			39428: outdata = 32'd26108;
			39429: outdata = 32'd26107;
			39430: outdata = 32'd26106;
			39431: outdata = 32'd26105;
			39432: outdata = 32'd26104;
			39433: outdata = 32'd26103;
			39434: outdata = 32'd26102;
			39435: outdata = 32'd26101;
			39436: outdata = 32'd26100;
			39437: outdata = 32'd26099;
			39438: outdata = 32'd26098;
			39439: outdata = 32'd26097;
			39440: outdata = 32'd26096;
			39441: outdata = 32'd26095;
			39442: outdata = 32'd26094;
			39443: outdata = 32'd26093;
			39444: outdata = 32'd26092;
			39445: outdata = 32'd26091;
			39446: outdata = 32'd26090;
			39447: outdata = 32'd26089;
			39448: outdata = 32'd26088;
			39449: outdata = 32'd26087;
			39450: outdata = 32'd26086;
			39451: outdata = 32'd26085;
			39452: outdata = 32'd26084;
			39453: outdata = 32'd26083;
			39454: outdata = 32'd26082;
			39455: outdata = 32'd26081;
			39456: outdata = 32'd26080;
			39457: outdata = 32'd26079;
			39458: outdata = 32'd26078;
			39459: outdata = 32'd26077;
			39460: outdata = 32'd26076;
			39461: outdata = 32'd26075;
			39462: outdata = 32'd26074;
			39463: outdata = 32'd26073;
			39464: outdata = 32'd26072;
			39465: outdata = 32'd26071;
			39466: outdata = 32'd26070;
			39467: outdata = 32'd26069;
			39468: outdata = 32'd26068;
			39469: outdata = 32'd26067;
			39470: outdata = 32'd26066;
			39471: outdata = 32'd26065;
			39472: outdata = 32'd26064;
			39473: outdata = 32'd26063;
			39474: outdata = 32'd26062;
			39475: outdata = 32'd26061;
			39476: outdata = 32'd26060;
			39477: outdata = 32'd26059;
			39478: outdata = 32'd26058;
			39479: outdata = 32'd26057;
			39480: outdata = 32'd26056;
			39481: outdata = 32'd26055;
			39482: outdata = 32'd26054;
			39483: outdata = 32'd26053;
			39484: outdata = 32'd26052;
			39485: outdata = 32'd26051;
			39486: outdata = 32'd26050;
			39487: outdata = 32'd26049;
			39488: outdata = 32'd26048;
			39489: outdata = 32'd26047;
			39490: outdata = 32'd26046;
			39491: outdata = 32'd26045;
			39492: outdata = 32'd26044;
			39493: outdata = 32'd26043;
			39494: outdata = 32'd26042;
			39495: outdata = 32'd26041;
			39496: outdata = 32'd26040;
			39497: outdata = 32'd26039;
			39498: outdata = 32'd26038;
			39499: outdata = 32'd26037;
			39500: outdata = 32'd26036;
			39501: outdata = 32'd26035;
			39502: outdata = 32'd26034;
			39503: outdata = 32'd26033;
			39504: outdata = 32'd26032;
			39505: outdata = 32'd26031;
			39506: outdata = 32'd26030;
			39507: outdata = 32'd26029;
			39508: outdata = 32'd26028;
			39509: outdata = 32'd26027;
			39510: outdata = 32'd26026;
			39511: outdata = 32'd26025;
			39512: outdata = 32'd26024;
			39513: outdata = 32'd26023;
			39514: outdata = 32'd26022;
			39515: outdata = 32'd26021;
			39516: outdata = 32'd26020;
			39517: outdata = 32'd26019;
			39518: outdata = 32'd26018;
			39519: outdata = 32'd26017;
			39520: outdata = 32'd26016;
			39521: outdata = 32'd26015;
			39522: outdata = 32'd26014;
			39523: outdata = 32'd26013;
			39524: outdata = 32'd26012;
			39525: outdata = 32'd26011;
			39526: outdata = 32'd26010;
			39527: outdata = 32'd26009;
			39528: outdata = 32'd26008;
			39529: outdata = 32'd26007;
			39530: outdata = 32'd26006;
			39531: outdata = 32'd26005;
			39532: outdata = 32'd26004;
			39533: outdata = 32'd26003;
			39534: outdata = 32'd26002;
			39535: outdata = 32'd26001;
			39536: outdata = 32'd26000;
			39537: outdata = 32'd25999;
			39538: outdata = 32'd25998;
			39539: outdata = 32'd25997;
			39540: outdata = 32'd25996;
			39541: outdata = 32'd25995;
			39542: outdata = 32'd25994;
			39543: outdata = 32'd25993;
			39544: outdata = 32'd25992;
			39545: outdata = 32'd25991;
			39546: outdata = 32'd25990;
			39547: outdata = 32'd25989;
			39548: outdata = 32'd25988;
			39549: outdata = 32'd25987;
			39550: outdata = 32'd25986;
			39551: outdata = 32'd25985;
			39552: outdata = 32'd25984;
			39553: outdata = 32'd25983;
			39554: outdata = 32'd25982;
			39555: outdata = 32'd25981;
			39556: outdata = 32'd25980;
			39557: outdata = 32'd25979;
			39558: outdata = 32'd25978;
			39559: outdata = 32'd25977;
			39560: outdata = 32'd25976;
			39561: outdata = 32'd25975;
			39562: outdata = 32'd25974;
			39563: outdata = 32'd25973;
			39564: outdata = 32'd25972;
			39565: outdata = 32'd25971;
			39566: outdata = 32'd25970;
			39567: outdata = 32'd25969;
			39568: outdata = 32'd25968;
			39569: outdata = 32'd25967;
			39570: outdata = 32'd25966;
			39571: outdata = 32'd25965;
			39572: outdata = 32'd25964;
			39573: outdata = 32'd25963;
			39574: outdata = 32'd25962;
			39575: outdata = 32'd25961;
			39576: outdata = 32'd25960;
			39577: outdata = 32'd25959;
			39578: outdata = 32'd25958;
			39579: outdata = 32'd25957;
			39580: outdata = 32'd25956;
			39581: outdata = 32'd25955;
			39582: outdata = 32'd25954;
			39583: outdata = 32'd25953;
			39584: outdata = 32'd25952;
			39585: outdata = 32'd25951;
			39586: outdata = 32'd25950;
			39587: outdata = 32'd25949;
			39588: outdata = 32'd25948;
			39589: outdata = 32'd25947;
			39590: outdata = 32'd25946;
			39591: outdata = 32'd25945;
			39592: outdata = 32'd25944;
			39593: outdata = 32'd25943;
			39594: outdata = 32'd25942;
			39595: outdata = 32'd25941;
			39596: outdata = 32'd25940;
			39597: outdata = 32'd25939;
			39598: outdata = 32'd25938;
			39599: outdata = 32'd25937;
			39600: outdata = 32'd25936;
			39601: outdata = 32'd25935;
			39602: outdata = 32'd25934;
			39603: outdata = 32'd25933;
			39604: outdata = 32'd25932;
			39605: outdata = 32'd25931;
			39606: outdata = 32'd25930;
			39607: outdata = 32'd25929;
			39608: outdata = 32'd25928;
			39609: outdata = 32'd25927;
			39610: outdata = 32'd25926;
			39611: outdata = 32'd25925;
			39612: outdata = 32'd25924;
			39613: outdata = 32'd25923;
			39614: outdata = 32'd25922;
			39615: outdata = 32'd25921;
			39616: outdata = 32'd25920;
			39617: outdata = 32'd25919;
			39618: outdata = 32'd25918;
			39619: outdata = 32'd25917;
			39620: outdata = 32'd25916;
			39621: outdata = 32'd25915;
			39622: outdata = 32'd25914;
			39623: outdata = 32'd25913;
			39624: outdata = 32'd25912;
			39625: outdata = 32'd25911;
			39626: outdata = 32'd25910;
			39627: outdata = 32'd25909;
			39628: outdata = 32'd25908;
			39629: outdata = 32'd25907;
			39630: outdata = 32'd25906;
			39631: outdata = 32'd25905;
			39632: outdata = 32'd25904;
			39633: outdata = 32'd25903;
			39634: outdata = 32'd25902;
			39635: outdata = 32'd25901;
			39636: outdata = 32'd25900;
			39637: outdata = 32'd25899;
			39638: outdata = 32'd25898;
			39639: outdata = 32'd25897;
			39640: outdata = 32'd25896;
			39641: outdata = 32'd25895;
			39642: outdata = 32'd25894;
			39643: outdata = 32'd25893;
			39644: outdata = 32'd25892;
			39645: outdata = 32'd25891;
			39646: outdata = 32'd25890;
			39647: outdata = 32'd25889;
			39648: outdata = 32'd25888;
			39649: outdata = 32'd25887;
			39650: outdata = 32'd25886;
			39651: outdata = 32'd25885;
			39652: outdata = 32'd25884;
			39653: outdata = 32'd25883;
			39654: outdata = 32'd25882;
			39655: outdata = 32'd25881;
			39656: outdata = 32'd25880;
			39657: outdata = 32'd25879;
			39658: outdata = 32'd25878;
			39659: outdata = 32'd25877;
			39660: outdata = 32'd25876;
			39661: outdata = 32'd25875;
			39662: outdata = 32'd25874;
			39663: outdata = 32'd25873;
			39664: outdata = 32'd25872;
			39665: outdata = 32'd25871;
			39666: outdata = 32'd25870;
			39667: outdata = 32'd25869;
			39668: outdata = 32'd25868;
			39669: outdata = 32'd25867;
			39670: outdata = 32'd25866;
			39671: outdata = 32'd25865;
			39672: outdata = 32'd25864;
			39673: outdata = 32'd25863;
			39674: outdata = 32'd25862;
			39675: outdata = 32'd25861;
			39676: outdata = 32'd25860;
			39677: outdata = 32'd25859;
			39678: outdata = 32'd25858;
			39679: outdata = 32'd25857;
			39680: outdata = 32'd25856;
			39681: outdata = 32'd25855;
			39682: outdata = 32'd25854;
			39683: outdata = 32'd25853;
			39684: outdata = 32'd25852;
			39685: outdata = 32'd25851;
			39686: outdata = 32'd25850;
			39687: outdata = 32'd25849;
			39688: outdata = 32'd25848;
			39689: outdata = 32'd25847;
			39690: outdata = 32'd25846;
			39691: outdata = 32'd25845;
			39692: outdata = 32'd25844;
			39693: outdata = 32'd25843;
			39694: outdata = 32'd25842;
			39695: outdata = 32'd25841;
			39696: outdata = 32'd25840;
			39697: outdata = 32'd25839;
			39698: outdata = 32'd25838;
			39699: outdata = 32'd25837;
			39700: outdata = 32'd25836;
			39701: outdata = 32'd25835;
			39702: outdata = 32'd25834;
			39703: outdata = 32'd25833;
			39704: outdata = 32'd25832;
			39705: outdata = 32'd25831;
			39706: outdata = 32'd25830;
			39707: outdata = 32'd25829;
			39708: outdata = 32'd25828;
			39709: outdata = 32'd25827;
			39710: outdata = 32'd25826;
			39711: outdata = 32'd25825;
			39712: outdata = 32'd25824;
			39713: outdata = 32'd25823;
			39714: outdata = 32'd25822;
			39715: outdata = 32'd25821;
			39716: outdata = 32'd25820;
			39717: outdata = 32'd25819;
			39718: outdata = 32'd25818;
			39719: outdata = 32'd25817;
			39720: outdata = 32'd25816;
			39721: outdata = 32'd25815;
			39722: outdata = 32'd25814;
			39723: outdata = 32'd25813;
			39724: outdata = 32'd25812;
			39725: outdata = 32'd25811;
			39726: outdata = 32'd25810;
			39727: outdata = 32'd25809;
			39728: outdata = 32'd25808;
			39729: outdata = 32'd25807;
			39730: outdata = 32'd25806;
			39731: outdata = 32'd25805;
			39732: outdata = 32'd25804;
			39733: outdata = 32'd25803;
			39734: outdata = 32'd25802;
			39735: outdata = 32'd25801;
			39736: outdata = 32'd25800;
			39737: outdata = 32'd25799;
			39738: outdata = 32'd25798;
			39739: outdata = 32'd25797;
			39740: outdata = 32'd25796;
			39741: outdata = 32'd25795;
			39742: outdata = 32'd25794;
			39743: outdata = 32'd25793;
			39744: outdata = 32'd25792;
			39745: outdata = 32'd25791;
			39746: outdata = 32'd25790;
			39747: outdata = 32'd25789;
			39748: outdata = 32'd25788;
			39749: outdata = 32'd25787;
			39750: outdata = 32'd25786;
			39751: outdata = 32'd25785;
			39752: outdata = 32'd25784;
			39753: outdata = 32'd25783;
			39754: outdata = 32'd25782;
			39755: outdata = 32'd25781;
			39756: outdata = 32'd25780;
			39757: outdata = 32'd25779;
			39758: outdata = 32'd25778;
			39759: outdata = 32'd25777;
			39760: outdata = 32'd25776;
			39761: outdata = 32'd25775;
			39762: outdata = 32'd25774;
			39763: outdata = 32'd25773;
			39764: outdata = 32'd25772;
			39765: outdata = 32'd25771;
			39766: outdata = 32'd25770;
			39767: outdata = 32'd25769;
			39768: outdata = 32'd25768;
			39769: outdata = 32'd25767;
			39770: outdata = 32'd25766;
			39771: outdata = 32'd25765;
			39772: outdata = 32'd25764;
			39773: outdata = 32'd25763;
			39774: outdata = 32'd25762;
			39775: outdata = 32'd25761;
			39776: outdata = 32'd25760;
			39777: outdata = 32'd25759;
			39778: outdata = 32'd25758;
			39779: outdata = 32'd25757;
			39780: outdata = 32'd25756;
			39781: outdata = 32'd25755;
			39782: outdata = 32'd25754;
			39783: outdata = 32'd25753;
			39784: outdata = 32'd25752;
			39785: outdata = 32'd25751;
			39786: outdata = 32'd25750;
			39787: outdata = 32'd25749;
			39788: outdata = 32'd25748;
			39789: outdata = 32'd25747;
			39790: outdata = 32'd25746;
			39791: outdata = 32'd25745;
			39792: outdata = 32'd25744;
			39793: outdata = 32'd25743;
			39794: outdata = 32'd25742;
			39795: outdata = 32'd25741;
			39796: outdata = 32'd25740;
			39797: outdata = 32'd25739;
			39798: outdata = 32'd25738;
			39799: outdata = 32'd25737;
			39800: outdata = 32'd25736;
			39801: outdata = 32'd25735;
			39802: outdata = 32'd25734;
			39803: outdata = 32'd25733;
			39804: outdata = 32'd25732;
			39805: outdata = 32'd25731;
			39806: outdata = 32'd25730;
			39807: outdata = 32'd25729;
			39808: outdata = 32'd25728;
			39809: outdata = 32'd25727;
			39810: outdata = 32'd25726;
			39811: outdata = 32'd25725;
			39812: outdata = 32'd25724;
			39813: outdata = 32'd25723;
			39814: outdata = 32'd25722;
			39815: outdata = 32'd25721;
			39816: outdata = 32'd25720;
			39817: outdata = 32'd25719;
			39818: outdata = 32'd25718;
			39819: outdata = 32'd25717;
			39820: outdata = 32'd25716;
			39821: outdata = 32'd25715;
			39822: outdata = 32'd25714;
			39823: outdata = 32'd25713;
			39824: outdata = 32'd25712;
			39825: outdata = 32'd25711;
			39826: outdata = 32'd25710;
			39827: outdata = 32'd25709;
			39828: outdata = 32'd25708;
			39829: outdata = 32'd25707;
			39830: outdata = 32'd25706;
			39831: outdata = 32'd25705;
			39832: outdata = 32'd25704;
			39833: outdata = 32'd25703;
			39834: outdata = 32'd25702;
			39835: outdata = 32'd25701;
			39836: outdata = 32'd25700;
			39837: outdata = 32'd25699;
			39838: outdata = 32'd25698;
			39839: outdata = 32'd25697;
			39840: outdata = 32'd25696;
			39841: outdata = 32'd25695;
			39842: outdata = 32'd25694;
			39843: outdata = 32'd25693;
			39844: outdata = 32'd25692;
			39845: outdata = 32'd25691;
			39846: outdata = 32'd25690;
			39847: outdata = 32'd25689;
			39848: outdata = 32'd25688;
			39849: outdata = 32'd25687;
			39850: outdata = 32'd25686;
			39851: outdata = 32'd25685;
			39852: outdata = 32'd25684;
			39853: outdata = 32'd25683;
			39854: outdata = 32'd25682;
			39855: outdata = 32'd25681;
			39856: outdata = 32'd25680;
			39857: outdata = 32'd25679;
			39858: outdata = 32'd25678;
			39859: outdata = 32'd25677;
			39860: outdata = 32'd25676;
			39861: outdata = 32'd25675;
			39862: outdata = 32'd25674;
			39863: outdata = 32'd25673;
			39864: outdata = 32'd25672;
			39865: outdata = 32'd25671;
			39866: outdata = 32'd25670;
			39867: outdata = 32'd25669;
			39868: outdata = 32'd25668;
			39869: outdata = 32'd25667;
			39870: outdata = 32'd25666;
			39871: outdata = 32'd25665;
			39872: outdata = 32'd25664;
			39873: outdata = 32'd25663;
			39874: outdata = 32'd25662;
			39875: outdata = 32'd25661;
			39876: outdata = 32'd25660;
			39877: outdata = 32'd25659;
			39878: outdata = 32'd25658;
			39879: outdata = 32'd25657;
			39880: outdata = 32'd25656;
			39881: outdata = 32'd25655;
			39882: outdata = 32'd25654;
			39883: outdata = 32'd25653;
			39884: outdata = 32'd25652;
			39885: outdata = 32'd25651;
			39886: outdata = 32'd25650;
			39887: outdata = 32'd25649;
			39888: outdata = 32'd25648;
			39889: outdata = 32'd25647;
			39890: outdata = 32'd25646;
			39891: outdata = 32'd25645;
			39892: outdata = 32'd25644;
			39893: outdata = 32'd25643;
			39894: outdata = 32'd25642;
			39895: outdata = 32'd25641;
			39896: outdata = 32'd25640;
			39897: outdata = 32'd25639;
			39898: outdata = 32'd25638;
			39899: outdata = 32'd25637;
			39900: outdata = 32'd25636;
			39901: outdata = 32'd25635;
			39902: outdata = 32'd25634;
			39903: outdata = 32'd25633;
			39904: outdata = 32'd25632;
			39905: outdata = 32'd25631;
			39906: outdata = 32'd25630;
			39907: outdata = 32'd25629;
			39908: outdata = 32'd25628;
			39909: outdata = 32'd25627;
			39910: outdata = 32'd25626;
			39911: outdata = 32'd25625;
			39912: outdata = 32'd25624;
			39913: outdata = 32'd25623;
			39914: outdata = 32'd25622;
			39915: outdata = 32'd25621;
			39916: outdata = 32'd25620;
			39917: outdata = 32'd25619;
			39918: outdata = 32'd25618;
			39919: outdata = 32'd25617;
			39920: outdata = 32'd25616;
			39921: outdata = 32'd25615;
			39922: outdata = 32'd25614;
			39923: outdata = 32'd25613;
			39924: outdata = 32'd25612;
			39925: outdata = 32'd25611;
			39926: outdata = 32'd25610;
			39927: outdata = 32'd25609;
			39928: outdata = 32'd25608;
			39929: outdata = 32'd25607;
			39930: outdata = 32'd25606;
			39931: outdata = 32'd25605;
			39932: outdata = 32'd25604;
			39933: outdata = 32'd25603;
			39934: outdata = 32'd25602;
			39935: outdata = 32'd25601;
			39936: outdata = 32'd25600;
			39937: outdata = 32'd25599;
			39938: outdata = 32'd25598;
			39939: outdata = 32'd25597;
			39940: outdata = 32'd25596;
			39941: outdata = 32'd25595;
			39942: outdata = 32'd25594;
			39943: outdata = 32'd25593;
			39944: outdata = 32'd25592;
			39945: outdata = 32'd25591;
			39946: outdata = 32'd25590;
			39947: outdata = 32'd25589;
			39948: outdata = 32'd25588;
			39949: outdata = 32'd25587;
			39950: outdata = 32'd25586;
			39951: outdata = 32'd25585;
			39952: outdata = 32'd25584;
			39953: outdata = 32'd25583;
			39954: outdata = 32'd25582;
			39955: outdata = 32'd25581;
			39956: outdata = 32'd25580;
			39957: outdata = 32'd25579;
			39958: outdata = 32'd25578;
			39959: outdata = 32'd25577;
			39960: outdata = 32'd25576;
			39961: outdata = 32'd25575;
			39962: outdata = 32'd25574;
			39963: outdata = 32'd25573;
			39964: outdata = 32'd25572;
			39965: outdata = 32'd25571;
			39966: outdata = 32'd25570;
			39967: outdata = 32'd25569;
			39968: outdata = 32'd25568;
			39969: outdata = 32'd25567;
			39970: outdata = 32'd25566;
			39971: outdata = 32'd25565;
			39972: outdata = 32'd25564;
			39973: outdata = 32'd25563;
			39974: outdata = 32'd25562;
			39975: outdata = 32'd25561;
			39976: outdata = 32'd25560;
			39977: outdata = 32'd25559;
			39978: outdata = 32'd25558;
			39979: outdata = 32'd25557;
			39980: outdata = 32'd25556;
			39981: outdata = 32'd25555;
			39982: outdata = 32'd25554;
			39983: outdata = 32'd25553;
			39984: outdata = 32'd25552;
			39985: outdata = 32'd25551;
			39986: outdata = 32'd25550;
			39987: outdata = 32'd25549;
			39988: outdata = 32'd25548;
			39989: outdata = 32'd25547;
			39990: outdata = 32'd25546;
			39991: outdata = 32'd25545;
			39992: outdata = 32'd25544;
			39993: outdata = 32'd25543;
			39994: outdata = 32'd25542;
			39995: outdata = 32'd25541;
			39996: outdata = 32'd25540;
			39997: outdata = 32'd25539;
			39998: outdata = 32'd25538;
			39999: outdata = 32'd25537;
			40000: outdata = 32'd25536;
			40001: outdata = 32'd25535;
			40002: outdata = 32'd25534;
			40003: outdata = 32'd25533;
			40004: outdata = 32'd25532;
			40005: outdata = 32'd25531;
			40006: outdata = 32'd25530;
			40007: outdata = 32'd25529;
			40008: outdata = 32'd25528;
			40009: outdata = 32'd25527;
			40010: outdata = 32'd25526;
			40011: outdata = 32'd25525;
			40012: outdata = 32'd25524;
			40013: outdata = 32'd25523;
			40014: outdata = 32'd25522;
			40015: outdata = 32'd25521;
			40016: outdata = 32'd25520;
			40017: outdata = 32'd25519;
			40018: outdata = 32'd25518;
			40019: outdata = 32'd25517;
			40020: outdata = 32'd25516;
			40021: outdata = 32'd25515;
			40022: outdata = 32'd25514;
			40023: outdata = 32'd25513;
			40024: outdata = 32'd25512;
			40025: outdata = 32'd25511;
			40026: outdata = 32'd25510;
			40027: outdata = 32'd25509;
			40028: outdata = 32'd25508;
			40029: outdata = 32'd25507;
			40030: outdata = 32'd25506;
			40031: outdata = 32'd25505;
			40032: outdata = 32'd25504;
			40033: outdata = 32'd25503;
			40034: outdata = 32'd25502;
			40035: outdata = 32'd25501;
			40036: outdata = 32'd25500;
			40037: outdata = 32'd25499;
			40038: outdata = 32'd25498;
			40039: outdata = 32'd25497;
			40040: outdata = 32'd25496;
			40041: outdata = 32'd25495;
			40042: outdata = 32'd25494;
			40043: outdata = 32'd25493;
			40044: outdata = 32'd25492;
			40045: outdata = 32'd25491;
			40046: outdata = 32'd25490;
			40047: outdata = 32'd25489;
			40048: outdata = 32'd25488;
			40049: outdata = 32'd25487;
			40050: outdata = 32'd25486;
			40051: outdata = 32'd25485;
			40052: outdata = 32'd25484;
			40053: outdata = 32'd25483;
			40054: outdata = 32'd25482;
			40055: outdata = 32'd25481;
			40056: outdata = 32'd25480;
			40057: outdata = 32'd25479;
			40058: outdata = 32'd25478;
			40059: outdata = 32'd25477;
			40060: outdata = 32'd25476;
			40061: outdata = 32'd25475;
			40062: outdata = 32'd25474;
			40063: outdata = 32'd25473;
			40064: outdata = 32'd25472;
			40065: outdata = 32'd25471;
			40066: outdata = 32'd25470;
			40067: outdata = 32'd25469;
			40068: outdata = 32'd25468;
			40069: outdata = 32'd25467;
			40070: outdata = 32'd25466;
			40071: outdata = 32'd25465;
			40072: outdata = 32'd25464;
			40073: outdata = 32'd25463;
			40074: outdata = 32'd25462;
			40075: outdata = 32'd25461;
			40076: outdata = 32'd25460;
			40077: outdata = 32'd25459;
			40078: outdata = 32'd25458;
			40079: outdata = 32'd25457;
			40080: outdata = 32'd25456;
			40081: outdata = 32'd25455;
			40082: outdata = 32'd25454;
			40083: outdata = 32'd25453;
			40084: outdata = 32'd25452;
			40085: outdata = 32'd25451;
			40086: outdata = 32'd25450;
			40087: outdata = 32'd25449;
			40088: outdata = 32'd25448;
			40089: outdata = 32'd25447;
			40090: outdata = 32'd25446;
			40091: outdata = 32'd25445;
			40092: outdata = 32'd25444;
			40093: outdata = 32'd25443;
			40094: outdata = 32'd25442;
			40095: outdata = 32'd25441;
			40096: outdata = 32'd25440;
			40097: outdata = 32'd25439;
			40098: outdata = 32'd25438;
			40099: outdata = 32'd25437;
			40100: outdata = 32'd25436;
			40101: outdata = 32'd25435;
			40102: outdata = 32'd25434;
			40103: outdata = 32'd25433;
			40104: outdata = 32'd25432;
			40105: outdata = 32'd25431;
			40106: outdata = 32'd25430;
			40107: outdata = 32'd25429;
			40108: outdata = 32'd25428;
			40109: outdata = 32'd25427;
			40110: outdata = 32'd25426;
			40111: outdata = 32'd25425;
			40112: outdata = 32'd25424;
			40113: outdata = 32'd25423;
			40114: outdata = 32'd25422;
			40115: outdata = 32'd25421;
			40116: outdata = 32'd25420;
			40117: outdata = 32'd25419;
			40118: outdata = 32'd25418;
			40119: outdata = 32'd25417;
			40120: outdata = 32'd25416;
			40121: outdata = 32'd25415;
			40122: outdata = 32'd25414;
			40123: outdata = 32'd25413;
			40124: outdata = 32'd25412;
			40125: outdata = 32'd25411;
			40126: outdata = 32'd25410;
			40127: outdata = 32'd25409;
			40128: outdata = 32'd25408;
			40129: outdata = 32'd25407;
			40130: outdata = 32'd25406;
			40131: outdata = 32'd25405;
			40132: outdata = 32'd25404;
			40133: outdata = 32'd25403;
			40134: outdata = 32'd25402;
			40135: outdata = 32'd25401;
			40136: outdata = 32'd25400;
			40137: outdata = 32'd25399;
			40138: outdata = 32'd25398;
			40139: outdata = 32'd25397;
			40140: outdata = 32'd25396;
			40141: outdata = 32'd25395;
			40142: outdata = 32'd25394;
			40143: outdata = 32'd25393;
			40144: outdata = 32'd25392;
			40145: outdata = 32'd25391;
			40146: outdata = 32'd25390;
			40147: outdata = 32'd25389;
			40148: outdata = 32'd25388;
			40149: outdata = 32'd25387;
			40150: outdata = 32'd25386;
			40151: outdata = 32'd25385;
			40152: outdata = 32'd25384;
			40153: outdata = 32'd25383;
			40154: outdata = 32'd25382;
			40155: outdata = 32'd25381;
			40156: outdata = 32'd25380;
			40157: outdata = 32'd25379;
			40158: outdata = 32'd25378;
			40159: outdata = 32'd25377;
			40160: outdata = 32'd25376;
			40161: outdata = 32'd25375;
			40162: outdata = 32'd25374;
			40163: outdata = 32'd25373;
			40164: outdata = 32'd25372;
			40165: outdata = 32'd25371;
			40166: outdata = 32'd25370;
			40167: outdata = 32'd25369;
			40168: outdata = 32'd25368;
			40169: outdata = 32'd25367;
			40170: outdata = 32'd25366;
			40171: outdata = 32'd25365;
			40172: outdata = 32'd25364;
			40173: outdata = 32'd25363;
			40174: outdata = 32'd25362;
			40175: outdata = 32'd25361;
			40176: outdata = 32'd25360;
			40177: outdata = 32'd25359;
			40178: outdata = 32'd25358;
			40179: outdata = 32'd25357;
			40180: outdata = 32'd25356;
			40181: outdata = 32'd25355;
			40182: outdata = 32'd25354;
			40183: outdata = 32'd25353;
			40184: outdata = 32'd25352;
			40185: outdata = 32'd25351;
			40186: outdata = 32'd25350;
			40187: outdata = 32'd25349;
			40188: outdata = 32'd25348;
			40189: outdata = 32'd25347;
			40190: outdata = 32'd25346;
			40191: outdata = 32'd25345;
			40192: outdata = 32'd25344;
			40193: outdata = 32'd25343;
			40194: outdata = 32'd25342;
			40195: outdata = 32'd25341;
			40196: outdata = 32'd25340;
			40197: outdata = 32'd25339;
			40198: outdata = 32'd25338;
			40199: outdata = 32'd25337;
			40200: outdata = 32'd25336;
			40201: outdata = 32'd25335;
			40202: outdata = 32'd25334;
			40203: outdata = 32'd25333;
			40204: outdata = 32'd25332;
			40205: outdata = 32'd25331;
			40206: outdata = 32'd25330;
			40207: outdata = 32'd25329;
			40208: outdata = 32'd25328;
			40209: outdata = 32'd25327;
			40210: outdata = 32'd25326;
			40211: outdata = 32'd25325;
			40212: outdata = 32'd25324;
			40213: outdata = 32'd25323;
			40214: outdata = 32'd25322;
			40215: outdata = 32'd25321;
			40216: outdata = 32'd25320;
			40217: outdata = 32'd25319;
			40218: outdata = 32'd25318;
			40219: outdata = 32'd25317;
			40220: outdata = 32'd25316;
			40221: outdata = 32'd25315;
			40222: outdata = 32'd25314;
			40223: outdata = 32'd25313;
			40224: outdata = 32'd25312;
			40225: outdata = 32'd25311;
			40226: outdata = 32'd25310;
			40227: outdata = 32'd25309;
			40228: outdata = 32'd25308;
			40229: outdata = 32'd25307;
			40230: outdata = 32'd25306;
			40231: outdata = 32'd25305;
			40232: outdata = 32'd25304;
			40233: outdata = 32'd25303;
			40234: outdata = 32'd25302;
			40235: outdata = 32'd25301;
			40236: outdata = 32'd25300;
			40237: outdata = 32'd25299;
			40238: outdata = 32'd25298;
			40239: outdata = 32'd25297;
			40240: outdata = 32'd25296;
			40241: outdata = 32'd25295;
			40242: outdata = 32'd25294;
			40243: outdata = 32'd25293;
			40244: outdata = 32'd25292;
			40245: outdata = 32'd25291;
			40246: outdata = 32'd25290;
			40247: outdata = 32'd25289;
			40248: outdata = 32'd25288;
			40249: outdata = 32'd25287;
			40250: outdata = 32'd25286;
			40251: outdata = 32'd25285;
			40252: outdata = 32'd25284;
			40253: outdata = 32'd25283;
			40254: outdata = 32'd25282;
			40255: outdata = 32'd25281;
			40256: outdata = 32'd25280;
			40257: outdata = 32'd25279;
			40258: outdata = 32'd25278;
			40259: outdata = 32'd25277;
			40260: outdata = 32'd25276;
			40261: outdata = 32'd25275;
			40262: outdata = 32'd25274;
			40263: outdata = 32'd25273;
			40264: outdata = 32'd25272;
			40265: outdata = 32'd25271;
			40266: outdata = 32'd25270;
			40267: outdata = 32'd25269;
			40268: outdata = 32'd25268;
			40269: outdata = 32'd25267;
			40270: outdata = 32'd25266;
			40271: outdata = 32'd25265;
			40272: outdata = 32'd25264;
			40273: outdata = 32'd25263;
			40274: outdata = 32'd25262;
			40275: outdata = 32'd25261;
			40276: outdata = 32'd25260;
			40277: outdata = 32'd25259;
			40278: outdata = 32'd25258;
			40279: outdata = 32'd25257;
			40280: outdata = 32'd25256;
			40281: outdata = 32'd25255;
			40282: outdata = 32'd25254;
			40283: outdata = 32'd25253;
			40284: outdata = 32'd25252;
			40285: outdata = 32'd25251;
			40286: outdata = 32'd25250;
			40287: outdata = 32'd25249;
			40288: outdata = 32'd25248;
			40289: outdata = 32'd25247;
			40290: outdata = 32'd25246;
			40291: outdata = 32'd25245;
			40292: outdata = 32'd25244;
			40293: outdata = 32'd25243;
			40294: outdata = 32'd25242;
			40295: outdata = 32'd25241;
			40296: outdata = 32'd25240;
			40297: outdata = 32'd25239;
			40298: outdata = 32'd25238;
			40299: outdata = 32'd25237;
			40300: outdata = 32'd25236;
			40301: outdata = 32'd25235;
			40302: outdata = 32'd25234;
			40303: outdata = 32'd25233;
			40304: outdata = 32'd25232;
			40305: outdata = 32'd25231;
			40306: outdata = 32'd25230;
			40307: outdata = 32'd25229;
			40308: outdata = 32'd25228;
			40309: outdata = 32'd25227;
			40310: outdata = 32'd25226;
			40311: outdata = 32'd25225;
			40312: outdata = 32'd25224;
			40313: outdata = 32'd25223;
			40314: outdata = 32'd25222;
			40315: outdata = 32'd25221;
			40316: outdata = 32'd25220;
			40317: outdata = 32'd25219;
			40318: outdata = 32'd25218;
			40319: outdata = 32'd25217;
			40320: outdata = 32'd25216;
			40321: outdata = 32'd25215;
			40322: outdata = 32'd25214;
			40323: outdata = 32'd25213;
			40324: outdata = 32'd25212;
			40325: outdata = 32'd25211;
			40326: outdata = 32'd25210;
			40327: outdata = 32'd25209;
			40328: outdata = 32'd25208;
			40329: outdata = 32'd25207;
			40330: outdata = 32'd25206;
			40331: outdata = 32'd25205;
			40332: outdata = 32'd25204;
			40333: outdata = 32'd25203;
			40334: outdata = 32'd25202;
			40335: outdata = 32'd25201;
			40336: outdata = 32'd25200;
			40337: outdata = 32'd25199;
			40338: outdata = 32'd25198;
			40339: outdata = 32'd25197;
			40340: outdata = 32'd25196;
			40341: outdata = 32'd25195;
			40342: outdata = 32'd25194;
			40343: outdata = 32'd25193;
			40344: outdata = 32'd25192;
			40345: outdata = 32'd25191;
			40346: outdata = 32'd25190;
			40347: outdata = 32'd25189;
			40348: outdata = 32'd25188;
			40349: outdata = 32'd25187;
			40350: outdata = 32'd25186;
			40351: outdata = 32'd25185;
			40352: outdata = 32'd25184;
			40353: outdata = 32'd25183;
			40354: outdata = 32'd25182;
			40355: outdata = 32'd25181;
			40356: outdata = 32'd25180;
			40357: outdata = 32'd25179;
			40358: outdata = 32'd25178;
			40359: outdata = 32'd25177;
			40360: outdata = 32'd25176;
			40361: outdata = 32'd25175;
			40362: outdata = 32'd25174;
			40363: outdata = 32'd25173;
			40364: outdata = 32'd25172;
			40365: outdata = 32'd25171;
			40366: outdata = 32'd25170;
			40367: outdata = 32'd25169;
			40368: outdata = 32'd25168;
			40369: outdata = 32'd25167;
			40370: outdata = 32'd25166;
			40371: outdata = 32'd25165;
			40372: outdata = 32'd25164;
			40373: outdata = 32'd25163;
			40374: outdata = 32'd25162;
			40375: outdata = 32'd25161;
			40376: outdata = 32'd25160;
			40377: outdata = 32'd25159;
			40378: outdata = 32'd25158;
			40379: outdata = 32'd25157;
			40380: outdata = 32'd25156;
			40381: outdata = 32'd25155;
			40382: outdata = 32'd25154;
			40383: outdata = 32'd25153;
			40384: outdata = 32'd25152;
			40385: outdata = 32'd25151;
			40386: outdata = 32'd25150;
			40387: outdata = 32'd25149;
			40388: outdata = 32'd25148;
			40389: outdata = 32'd25147;
			40390: outdata = 32'd25146;
			40391: outdata = 32'd25145;
			40392: outdata = 32'd25144;
			40393: outdata = 32'd25143;
			40394: outdata = 32'd25142;
			40395: outdata = 32'd25141;
			40396: outdata = 32'd25140;
			40397: outdata = 32'd25139;
			40398: outdata = 32'd25138;
			40399: outdata = 32'd25137;
			40400: outdata = 32'd25136;
			40401: outdata = 32'd25135;
			40402: outdata = 32'd25134;
			40403: outdata = 32'd25133;
			40404: outdata = 32'd25132;
			40405: outdata = 32'd25131;
			40406: outdata = 32'd25130;
			40407: outdata = 32'd25129;
			40408: outdata = 32'd25128;
			40409: outdata = 32'd25127;
			40410: outdata = 32'd25126;
			40411: outdata = 32'd25125;
			40412: outdata = 32'd25124;
			40413: outdata = 32'd25123;
			40414: outdata = 32'd25122;
			40415: outdata = 32'd25121;
			40416: outdata = 32'd25120;
			40417: outdata = 32'd25119;
			40418: outdata = 32'd25118;
			40419: outdata = 32'd25117;
			40420: outdata = 32'd25116;
			40421: outdata = 32'd25115;
			40422: outdata = 32'd25114;
			40423: outdata = 32'd25113;
			40424: outdata = 32'd25112;
			40425: outdata = 32'd25111;
			40426: outdata = 32'd25110;
			40427: outdata = 32'd25109;
			40428: outdata = 32'd25108;
			40429: outdata = 32'd25107;
			40430: outdata = 32'd25106;
			40431: outdata = 32'd25105;
			40432: outdata = 32'd25104;
			40433: outdata = 32'd25103;
			40434: outdata = 32'd25102;
			40435: outdata = 32'd25101;
			40436: outdata = 32'd25100;
			40437: outdata = 32'd25099;
			40438: outdata = 32'd25098;
			40439: outdata = 32'd25097;
			40440: outdata = 32'd25096;
			40441: outdata = 32'd25095;
			40442: outdata = 32'd25094;
			40443: outdata = 32'd25093;
			40444: outdata = 32'd25092;
			40445: outdata = 32'd25091;
			40446: outdata = 32'd25090;
			40447: outdata = 32'd25089;
			40448: outdata = 32'd25088;
			40449: outdata = 32'd25087;
			40450: outdata = 32'd25086;
			40451: outdata = 32'd25085;
			40452: outdata = 32'd25084;
			40453: outdata = 32'd25083;
			40454: outdata = 32'd25082;
			40455: outdata = 32'd25081;
			40456: outdata = 32'd25080;
			40457: outdata = 32'd25079;
			40458: outdata = 32'd25078;
			40459: outdata = 32'd25077;
			40460: outdata = 32'd25076;
			40461: outdata = 32'd25075;
			40462: outdata = 32'd25074;
			40463: outdata = 32'd25073;
			40464: outdata = 32'd25072;
			40465: outdata = 32'd25071;
			40466: outdata = 32'd25070;
			40467: outdata = 32'd25069;
			40468: outdata = 32'd25068;
			40469: outdata = 32'd25067;
			40470: outdata = 32'd25066;
			40471: outdata = 32'd25065;
			40472: outdata = 32'd25064;
			40473: outdata = 32'd25063;
			40474: outdata = 32'd25062;
			40475: outdata = 32'd25061;
			40476: outdata = 32'd25060;
			40477: outdata = 32'd25059;
			40478: outdata = 32'd25058;
			40479: outdata = 32'd25057;
			40480: outdata = 32'd25056;
			40481: outdata = 32'd25055;
			40482: outdata = 32'd25054;
			40483: outdata = 32'd25053;
			40484: outdata = 32'd25052;
			40485: outdata = 32'd25051;
			40486: outdata = 32'd25050;
			40487: outdata = 32'd25049;
			40488: outdata = 32'd25048;
			40489: outdata = 32'd25047;
			40490: outdata = 32'd25046;
			40491: outdata = 32'd25045;
			40492: outdata = 32'd25044;
			40493: outdata = 32'd25043;
			40494: outdata = 32'd25042;
			40495: outdata = 32'd25041;
			40496: outdata = 32'd25040;
			40497: outdata = 32'd25039;
			40498: outdata = 32'd25038;
			40499: outdata = 32'd25037;
			40500: outdata = 32'd25036;
			40501: outdata = 32'd25035;
			40502: outdata = 32'd25034;
			40503: outdata = 32'd25033;
			40504: outdata = 32'd25032;
			40505: outdata = 32'd25031;
			40506: outdata = 32'd25030;
			40507: outdata = 32'd25029;
			40508: outdata = 32'd25028;
			40509: outdata = 32'd25027;
			40510: outdata = 32'd25026;
			40511: outdata = 32'd25025;
			40512: outdata = 32'd25024;
			40513: outdata = 32'd25023;
			40514: outdata = 32'd25022;
			40515: outdata = 32'd25021;
			40516: outdata = 32'd25020;
			40517: outdata = 32'd25019;
			40518: outdata = 32'd25018;
			40519: outdata = 32'd25017;
			40520: outdata = 32'd25016;
			40521: outdata = 32'd25015;
			40522: outdata = 32'd25014;
			40523: outdata = 32'd25013;
			40524: outdata = 32'd25012;
			40525: outdata = 32'd25011;
			40526: outdata = 32'd25010;
			40527: outdata = 32'd25009;
			40528: outdata = 32'd25008;
			40529: outdata = 32'd25007;
			40530: outdata = 32'd25006;
			40531: outdata = 32'd25005;
			40532: outdata = 32'd25004;
			40533: outdata = 32'd25003;
			40534: outdata = 32'd25002;
			40535: outdata = 32'd25001;
			40536: outdata = 32'd25000;
			40537: outdata = 32'd24999;
			40538: outdata = 32'd24998;
			40539: outdata = 32'd24997;
			40540: outdata = 32'd24996;
			40541: outdata = 32'd24995;
			40542: outdata = 32'd24994;
			40543: outdata = 32'd24993;
			40544: outdata = 32'd24992;
			40545: outdata = 32'd24991;
			40546: outdata = 32'd24990;
			40547: outdata = 32'd24989;
			40548: outdata = 32'd24988;
			40549: outdata = 32'd24987;
			40550: outdata = 32'd24986;
			40551: outdata = 32'd24985;
			40552: outdata = 32'd24984;
			40553: outdata = 32'd24983;
			40554: outdata = 32'd24982;
			40555: outdata = 32'd24981;
			40556: outdata = 32'd24980;
			40557: outdata = 32'd24979;
			40558: outdata = 32'd24978;
			40559: outdata = 32'd24977;
			40560: outdata = 32'd24976;
			40561: outdata = 32'd24975;
			40562: outdata = 32'd24974;
			40563: outdata = 32'd24973;
			40564: outdata = 32'd24972;
			40565: outdata = 32'd24971;
			40566: outdata = 32'd24970;
			40567: outdata = 32'd24969;
			40568: outdata = 32'd24968;
			40569: outdata = 32'd24967;
			40570: outdata = 32'd24966;
			40571: outdata = 32'd24965;
			40572: outdata = 32'd24964;
			40573: outdata = 32'd24963;
			40574: outdata = 32'd24962;
			40575: outdata = 32'd24961;
			40576: outdata = 32'd24960;
			40577: outdata = 32'd24959;
			40578: outdata = 32'd24958;
			40579: outdata = 32'd24957;
			40580: outdata = 32'd24956;
			40581: outdata = 32'd24955;
			40582: outdata = 32'd24954;
			40583: outdata = 32'd24953;
			40584: outdata = 32'd24952;
			40585: outdata = 32'd24951;
			40586: outdata = 32'd24950;
			40587: outdata = 32'd24949;
			40588: outdata = 32'd24948;
			40589: outdata = 32'd24947;
			40590: outdata = 32'd24946;
			40591: outdata = 32'd24945;
			40592: outdata = 32'd24944;
			40593: outdata = 32'd24943;
			40594: outdata = 32'd24942;
			40595: outdata = 32'd24941;
			40596: outdata = 32'd24940;
			40597: outdata = 32'd24939;
			40598: outdata = 32'd24938;
			40599: outdata = 32'd24937;
			40600: outdata = 32'd24936;
			40601: outdata = 32'd24935;
			40602: outdata = 32'd24934;
			40603: outdata = 32'd24933;
			40604: outdata = 32'd24932;
			40605: outdata = 32'd24931;
			40606: outdata = 32'd24930;
			40607: outdata = 32'd24929;
			40608: outdata = 32'd24928;
			40609: outdata = 32'd24927;
			40610: outdata = 32'd24926;
			40611: outdata = 32'd24925;
			40612: outdata = 32'd24924;
			40613: outdata = 32'd24923;
			40614: outdata = 32'd24922;
			40615: outdata = 32'd24921;
			40616: outdata = 32'd24920;
			40617: outdata = 32'd24919;
			40618: outdata = 32'd24918;
			40619: outdata = 32'd24917;
			40620: outdata = 32'd24916;
			40621: outdata = 32'd24915;
			40622: outdata = 32'd24914;
			40623: outdata = 32'd24913;
			40624: outdata = 32'd24912;
			40625: outdata = 32'd24911;
			40626: outdata = 32'd24910;
			40627: outdata = 32'd24909;
			40628: outdata = 32'd24908;
			40629: outdata = 32'd24907;
			40630: outdata = 32'd24906;
			40631: outdata = 32'd24905;
			40632: outdata = 32'd24904;
			40633: outdata = 32'd24903;
			40634: outdata = 32'd24902;
			40635: outdata = 32'd24901;
			40636: outdata = 32'd24900;
			40637: outdata = 32'd24899;
			40638: outdata = 32'd24898;
			40639: outdata = 32'd24897;
			40640: outdata = 32'd24896;
			40641: outdata = 32'd24895;
			40642: outdata = 32'd24894;
			40643: outdata = 32'd24893;
			40644: outdata = 32'd24892;
			40645: outdata = 32'd24891;
			40646: outdata = 32'd24890;
			40647: outdata = 32'd24889;
			40648: outdata = 32'd24888;
			40649: outdata = 32'd24887;
			40650: outdata = 32'd24886;
			40651: outdata = 32'd24885;
			40652: outdata = 32'd24884;
			40653: outdata = 32'd24883;
			40654: outdata = 32'd24882;
			40655: outdata = 32'd24881;
			40656: outdata = 32'd24880;
			40657: outdata = 32'd24879;
			40658: outdata = 32'd24878;
			40659: outdata = 32'd24877;
			40660: outdata = 32'd24876;
			40661: outdata = 32'd24875;
			40662: outdata = 32'd24874;
			40663: outdata = 32'd24873;
			40664: outdata = 32'd24872;
			40665: outdata = 32'd24871;
			40666: outdata = 32'd24870;
			40667: outdata = 32'd24869;
			40668: outdata = 32'd24868;
			40669: outdata = 32'd24867;
			40670: outdata = 32'd24866;
			40671: outdata = 32'd24865;
			40672: outdata = 32'd24864;
			40673: outdata = 32'd24863;
			40674: outdata = 32'd24862;
			40675: outdata = 32'd24861;
			40676: outdata = 32'd24860;
			40677: outdata = 32'd24859;
			40678: outdata = 32'd24858;
			40679: outdata = 32'd24857;
			40680: outdata = 32'd24856;
			40681: outdata = 32'd24855;
			40682: outdata = 32'd24854;
			40683: outdata = 32'd24853;
			40684: outdata = 32'd24852;
			40685: outdata = 32'd24851;
			40686: outdata = 32'd24850;
			40687: outdata = 32'd24849;
			40688: outdata = 32'd24848;
			40689: outdata = 32'd24847;
			40690: outdata = 32'd24846;
			40691: outdata = 32'd24845;
			40692: outdata = 32'd24844;
			40693: outdata = 32'd24843;
			40694: outdata = 32'd24842;
			40695: outdata = 32'd24841;
			40696: outdata = 32'd24840;
			40697: outdata = 32'd24839;
			40698: outdata = 32'd24838;
			40699: outdata = 32'd24837;
			40700: outdata = 32'd24836;
			40701: outdata = 32'd24835;
			40702: outdata = 32'd24834;
			40703: outdata = 32'd24833;
			40704: outdata = 32'd24832;
			40705: outdata = 32'd24831;
			40706: outdata = 32'd24830;
			40707: outdata = 32'd24829;
			40708: outdata = 32'd24828;
			40709: outdata = 32'd24827;
			40710: outdata = 32'd24826;
			40711: outdata = 32'd24825;
			40712: outdata = 32'd24824;
			40713: outdata = 32'd24823;
			40714: outdata = 32'd24822;
			40715: outdata = 32'd24821;
			40716: outdata = 32'd24820;
			40717: outdata = 32'd24819;
			40718: outdata = 32'd24818;
			40719: outdata = 32'd24817;
			40720: outdata = 32'd24816;
			40721: outdata = 32'd24815;
			40722: outdata = 32'd24814;
			40723: outdata = 32'd24813;
			40724: outdata = 32'd24812;
			40725: outdata = 32'd24811;
			40726: outdata = 32'd24810;
			40727: outdata = 32'd24809;
			40728: outdata = 32'd24808;
			40729: outdata = 32'd24807;
			40730: outdata = 32'd24806;
			40731: outdata = 32'd24805;
			40732: outdata = 32'd24804;
			40733: outdata = 32'd24803;
			40734: outdata = 32'd24802;
			40735: outdata = 32'd24801;
			40736: outdata = 32'd24800;
			40737: outdata = 32'd24799;
			40738: outdata = 32'd24798;
			40739: outdata = 32'd24797;
			40740: outdata = 32'd24796;
			40741: outdata = 32'd24795;
			40742: outdata = 32'd24794;
			40743: outdata = 32'd24793;
			40744: outdata = 32'd24792;
			40745: outdata = 32'd24791;
			40746: outdata = 32'd24790;
			40747: outdata = 32'd24789;
			40748: outdata = 32'd24788;
			40749: outdata = 32'd24787;
			40750: outdata = 32'd24786;
			40751: outdata = 32'd24785;
			40752: outdata = 32'd24784;
			40753: outdata = 32'd24783;
			40754: outdata = 32'd24782;
			40755: outdata = 32'd24781;
			40756: outdata = 32'd24780;
			40757: outdata = 32'd24779;
			40758: outdata = 32'd24778;
			40759: outdata = 32'd24777;
			40760: outdata = 32'd24776;
			40761: outdata = 32'd24775;
			40762: outdata = 32'd24774;
			40763: outdata = 32'd24773;
			40764: outdata = 32'd24772;
			40765: outdata = 32'd24771;
			40766: outdata = 32'd24770;
			40767: outdata = 32'd24769;
			40768: outdata = 32'd24768;
			40769: outdata = 32'd24767;
			40770: outdata = 32'd24766;
			40771: outdata = 32'd24765;
			40772: outdata = 32'd24764;
			40773: outdata = 32'd24763;
			40774: outdata = 32'd24762;
			40775: outdata = 32'd24761;
			40776: outdata = 32'd24760;
			40777: outdata = 32'd24759;
			40778: outdata = 32'd24758;
			40779: outdata = 32'd24757;
			40780: outdata = 32'd24756;
			40781: outdata = 32'd24755;
			40782: outdata = 32'd24754;
			40783: outdata = 32'd24753;
			40784: outdata = 32'd24752;
			40785: outdata = 32'd24751;
			40786: outdata = 32'd24750;
			40787: outdata = 32'd24749;
			40788: outdata = 32'd24748;
			40789: outdata = 32'd24747;
			40790: outdata = 32'd24746;
			40791: outdata = 32'd24745;
			40792: outdata = 32'd24744;
			40793: outdata = 32'd24743;
			40794: outdata = 32'd24742;
			40795: outdata = 32'd24741;
			40796: outdata = 32'd24740;
			40797: outdata = 32'd24739;
			40798: outdata = 32'd24738;
			40799: outdata = 32'd24737;
			40800: outdata = 32'd24736;
			40801: outdata = 32'd24735;
			40802: outdata = 32'd24734;
			40803: outdata = 32'd24733;
			40804: outdata = 32'd24732;
			40805: outdata = 32'd24731;
			40806: outdata = 32'd24730;
			40807: outdata = 32'd24729;
			40808: outdata = 32'd24728;
			40809: outdata = 32'd24727;
			40810: outdata = 32'd24726;
			40811: outdata = 32'd24725;
			40812: outdata = 32'd24724;
			40813: outdata = 32'd24723;
			40814: outdata = 32'd24722;
			40815: outdata = 32'd24721;
			40816: outdata = 32'd24720;
			40817: outdata = 32'd24719;
			40818: outdata = 32'd24718;
			40819: outdata = 32'd24717;
			40820: outdata = 32'd24716;
			40821: outdata = 32'd24715;
			40822: outdata = 32'd24714;
			40823: outdata = 32'd24713;
			40824: outdata = 32'd24712;
			40825: outdata = 32'd24711;
			40826: outdata = 32'd24710;
			40827: outdata = 32'd24709;
			40828: outdata = 32'd24708;
			40829: outdata = 32'd24707;
			40830: outdata = 32'd24706;
			40831: outdata = 32'd24705;
			40832: outdata = 32'd24704;
			40833: outdata = 32'd24703;
			40834: outdata = 32'd24702;
			40835: outdata = 32'd24701;
			40836: outdata = 32'd24700;
			40837: outdata = 32'd24699;
			40838: outdata = 32'd24698;
			40839: outdata = 32'd24697;
			40840: outdata = 32'd24696;
			40841: outdata = 32'd24695;
			40842: outdata = 32'd24694;
			40843: outdata = 32'd24693;
			40844: outdata = 32'd24692;
			40845: outdata = 32'd24691;
			40846: outdata = 32'd24690;
			40847: outdata = 32'd24689;
			40848: outdata = 32'd24688;
			40849: outdata = 32'd24687;
			40850: outdata = 32'd24686;
			40851: outdata = 32'd24685;
			40852: outdata = 32'd24684;
			40853: outdata = 32'd24683;
			40854: outdata = 32'd24682;
			40855: outdata = 32'd24681;
			40856: outdata = 32'd24680;
			40857: outdata = 32'd24679;
			40858: outdata = 32'd24678;
			40859: outdata = 32'd24677;
			40860: outdata = 32'd24676;
			40861: outdata = 32'd24675;
			40862: outdata = 32'd24674;
			40863: outdata = 32'd24673;
			40864: outdata = 32'd24672;
			40865: outdata = 32'd24671;
			40866: outdata = 32'd24670;
			40867: outdata = 32'd24669;
			40868: outdata = 32'd24668;
			40869: outdata = 32'd24667;
			40870: outdata = 32'd24666;
			40871: outdata = 32'd24665;
			40872: outdata = 32'd24664;
			40873: outdata = 32'd24663;
			40874: outdata = 32'd24662;
			40875: outdata = 32'd24661;
			40876: outdata = 32'd24660;
			40877: outdata = 32'd24659;
			40878: outdata = 32'd24658;
			40879: outdata = 32'd24657;
			40880: outdata = 32'd24656;
			40881: outdata = 32'd24655;
			40882: outdata = 32'd24654;
			40883: outdata = 32'd24653;
			40884: outdata = 32'd24652;
			40885: outdata = 32'd24651;
			40886: outdata = 32'd24650;
			40887: outdata = 32'd24649;
			40888: outdata = 32'd24648;
			40889: outdata = 32'd24647;
			40890: outdata = 32'd24646;
			40891: outdata = 32'd24645;
			40892: outdata = 32'd24644;
			40893: outdata = 32'd24643;
			40894: outdata = 32'd24642;
			40895: outdata = 32'd24641;
			40896: outdata = 32'd24640;
			40897: outdata = 32'd24639;
			40898: outdata = 32'd24638;
			40899: outdata = 32'd24637;
			40900: outdata = 32'd24636;
			40901: outdata = 32'd24635;
			40902: outdata = 32'd24634;
			40903: outdata = 32'd24633;
			40904: outdata = 32'd24632;
			40905: outdata = 32'd24631;
			40906: outdata = 32'd24630;
			40907: outdata = 32'd24629;
			40908: outdata = 32'd24628;
			40909: outdata = 32'd24627;
			40910: outdata = 32'd24626;
			40911: outdata = 32'd24625;
			40912: outdata = 32'd24624;
			40913: outdata = 32'd24623;
			40914: outdata = 32'd24622;
			40915: outdata = 32'd24621;
			40916: outdata = 32'd24620;
			40917: outdata = 32'd24619;
			40918: outdata = 32'd24618;
			40919: outdata = 32'd24617;
			40920: outdata = 32'd24616;
			40921: outdata = 32'd24615;
			40922: outdata = 32'd24614;
			40923: outdata = 32'd24613;
			40924: outdata = 32'd24612;
			40925: outdata = 32'd24611;
			40926: outdata = 32'd24610;
			40927: outdata = 32'd24609;
			40928: outdata = 32'd24608;
			40929: outdata = 32'd24607;
			40930: outdata = 32'd24606;
			40931: outdata = 32'd24605;
			40932: outdata = 32'd24604;
			40933: outdata = 32'd24603;
			40934: outdata = 32'd24602;
			40935: outdata = 32'd24601;
			40936: outdata = 32'd24600;
			40937: outdata = 32'd24599;
			40938: outdata = 32'd24598;
			40939: outdata = 32'd24597;
			40940: outdata = 32'd24596;
			40941: outdata = 32'd24595;
			40942: outdata = 32'd24594;
			40943: outdata = 32'd24593;
			40944: outdata = 32'd24592;
			40945: outdata = 32'd24591;
			40946: outdata = 32'd24590;
			40947: outdata = 32'd24589;
			40948: outdata = 32'd24588;
			40949: outdata = 32'd24587;
			40950: outdata = 32'd24586;
			40951: outdata = 32'd24585;
			40952: outdata = 32'd24584;
			40953: outdata = 32'd24583;
			40954: outdata = 32'd24582;
			40955: outdata = 32'd24581;
			40956: outdata = 32'd24580;
			40957: outdata = 32'd24579;
			40958: outdata = 32'd24578;
			40959: outdata = 32'd24577;
			40960: outdata = 32'd24576;
			40961: outdata = 32'd24575;
			40962: outdata = 32'd24574;
			40963: outdata = 32'd24573;
			40964: outdata = 32'd24572;
			40965: outdata = 32'd24571;
			40966: outdata = 32'd24570;
			40967: outdata = 32'd24569;
			40968: outdata = 32'd24568;
			40969: outdata = 32'd24567;
			40970: outdata = 32'd24566;
			40971: outdata = 32'd24565;
			40972: outdata = 32'd24564;
			40973: outdata = 32'd24563;
			40974: outdata = 32'd24562;
			40975: outdata = 32'd24561;
			40976: outdata = 32'd24560;
			40977: outdata = 32'd24559;
			40978: outdata = 32'd24558;
			40979: outdata = 32'd24557;
			40980: outdata = 32'd24556;
			40981: outdata = 32'd24555;
			40982: outdata = 32'd24554;
			40983: outdata = 32'd24553;
			40984: outdata = 32'd24552;
			40985: outdata = 32'd24551;
			40986: outdata = 32'd24550;
			40987: outdata = 32'd24549;
			40988: outdata = 32'd24548;
			40989: outdata = 32'd24547;
			40990: outdata = 32'd24546;
			40991: outdata = 32'd24545;
			40992: outdata = 32'd24544;
			40993: outdata = 32'd24543;
			40994: outdata = 32'd24542;
			40995: outdata = 32'd24541;
			40996: outdata = 32'd24540;
			40997: outdata = 32'd24539;
			40998: outdata = 32'd24538;
			40999: outdata = 32'd24537;
			41000: outdata = 32'd24536;
			41001: outdata = 32'd24535;
			41002: outdata = 32'd24534;
			41003: outdata = 32'd24533;
			41004: outdata = 32'd24532;
			41005: outdata = 32'd24531;
			41006: outdata = 32'd24530;
			41007: outdata = 32'd24529;
			41008: outdata = 32'd24528;
			41009: outdata = 32'd24527;
			41010: outdata = 32'd24526;
			41011: outdata = 32'd24525;
			41012: outdata = 32'd24524;
			41013: outdata = 32'd24523;
			41014: outdata = 32'd24522;
			41015: outdata = 32'd24521;
			41016: outdata = 32'd24520;
			41017: outdata = 32'd24519;
			41018: outdata = 32'd24518;
			41019: outdata = 32'd24517;
			41020: outdata = 32'd24516;
			41021: outdata = 32'd24515;
			41022: outdata = 32'd24514;
			41023: outdata = 32'd24513;
			41024: outdata = 32'd24512;
			41025: outdata = 32'd24511;
			41026: outdata = 32'd24510;
			41027: outdata = 32'd24509;
			41028: outdata = 32'd24508;
			41029: outdata = 32'd24507;
			41030: outdata = 32'd24506;
			41031: outdata = 32'd24505;
			41032: outdata = 32'd24504;
			41033: outdata = 32'd24503;
			41034: outdata = 32'd24502;
			41035: outdata = 32'd24501;
			41036: outdata = 32'd24500;
			41037: outdata = 32'd24499;
			41038: outdata = 32'd24498;
			41039: outdata = 32'd24497;
			41040: outdata = 32'd24496;
			41041: outdata = 32'd24495;
			41042: outdata = 32'd24494;
			41043: outdata = 32'd24493;
			41044: outdata = 32'd24492;
			41045: outdata = 32'd24491;
			41046: outdata = 32'd24490;
			41047: outdata = 32'd24489;
			41048: outdata = 32'd24488;
			41049: outdata = 32'd24487;
			41050: outdata = 32'd24486;
			41051: outdata = 32'd24485;
			41052: outdata = 32'd24484;
			41053: outdata = 32'd24483;
			41054: outdata = 32'd24482;
			41055: outdata = 32'd24481;
			41056: outdata = 32'd24480;
			41057: outdata = 32'd24479;
			41058: outdata = 32'd24478;
			41059: outdata = 32'd24477;
			41060: outdata = 32'd24476;
			41061: outdata = 32'd24475;
			41062: outdata = 32'd24474;
			41063: outdata = 32'd24473;
			41064: outdata = 32'd24472;
			41065: outdata = 32'd24471;
			41066: outdata = 32'd24470;
			41067: outdata = 32'd24469;
			41068: outdata = 32'd24468;
			41069: outdata = 32'd24467;
			41070: outdata = 32'd24466;
			41071: outdata = 32'd24465;
			41072: outdata = 32'd24464;
			41073: outdata = 32'd24463;
			41074: outdata = 32'd24462;
			41075: outdata = 32'd24461;
			41076: outdata = 32'd24460;
			41077: outdata = 32'd24459;
			41078: outdata = 32'd24458;
			41079: outdata = 32'd24457;
			41080: outdata = 32'd24456;
			41081: outdata = 32'd24455;
			41082: outdata = 32'd24454;
			41083: outdata = 32'd24453;
			41084: outdata = 32'd24452;
			41085: outdata = 32'd24451;
			41086: outdata = 32'd24450;
			41087: outdata = 32'd24449;
			41088: outdata = 32'd24448;
			41089: outdata = 32'd24447;
			41090: outdata = 32'd24446;
			41091: outdata = 32'd24445;
			41092: outdata = 32'd24444;
			41093: outdata = 32'd24443;
			41094: outdata = 32'd24442;
			41095: outdata = 32'd24441;
			41096: outdata = 32'd24440;
			41097: outdata = 32'd24439;
			41098: outdata = 32'd24438;
			41099: outdata = 32'd24437;
			41100: outdata = 32'd24436;
			41101: outdata = 32'd24435;
			41102: outdata = 32'd24434;
			41103: outdata = 32'd24433;
			41104: outdata = 32'd24432;
			41105: outdata = 32'd24431;
			41106: outdata = 32'd24430;
			41107: outdata = 32'd24429;
			41108: outdata = 32'd24428;
			41109: outdata = 32'd24427;
			41110: outdata = 32'd24426;
			41111: outdata = 32'd24425;
			41112: outdata = 32'd24424;
			41113: outdata = 32'd24423;
			41114: outdata = 32'd24422;
			41115: outdata = 32'd24421;
			41116: outdata = 32'd24420;
			41117: outdata = 32'd24419;
			41118: outdata = 32'd24418;
			41119: outdata = 32'd24417;
			41120: outdata = 32'd24416;
			41121: outdata = 32'd24415;
			41122: outdata = 32'd24414;
			41123: outdata = 32'd24413;
			41124: outdata = 32'd24412;
			41125: outdata = 32'd24411;
			41126: outdata = 32'd24410;
			41127: outdata = 32'd24409;
			41128: outdata = 32'd24408;
			41129: outdata = 32'd24407;
			41130: outdata = 32'd24406;
			41131: outdata = 32'd24405;
			41132: outdata = 32'd24404;
			41133: outdata = 32'd24403;
			41134: outdata = 32'd24402;
			41135: outdata = 32'd24401;
			41136: outdata = 32'd24400;
			41137: outdata = 32'd24399;
			41138: outdata = 32'd24398;
			41139: outdata = 32'd24397;
			41140: outdata = 32'd24396;
			41141: outdata = 32'd24395;
			41142: outdata = 32'd24394;
			41143: outdata = 32'd24393;
			41144: outdata = 32'd24392;
			41145: outdata = 32'd24391;
			41146: outdata = 32'd24390;
			41147: outdata = 32'd24389;
			41148: outdata = 32'd24388;
			41149: outdata = 32'd24387;
			41150: outdata = 32'd24386;
			41151: outdata = 32'd24385;
			41152: outdata = 32'd24384;
			41153: outdata = 32'd24383;
			41154: outdata = 32'd24382;
			41155: outdata = 32'd24381;
			41156: outdata = 32'd24380;
			41157: outdata = 32'd24379;
			41158: outdata = 32'd24378;
			41159: outdata = 32'd24377;
			41160: outdata = 32'd24376;
			41161: outdata = 32'd24375;
			41162: outdata = 32'd24374;
			41163: outdata = 32'd24373;
			41164: outdata = 32'd24372;
			41165: outdata = 32'd24371;
			41166: outdata = 32'd24370;
			41167: outdata = 32'd24369;
			41168: outdata = 32'd24368;
			41169: outdata = 32'd24367;
			41170: outdata = 32'd24366;
			41171: outdata = 32'd24365;
			41172: outdata = 32'd24364;
			41173: outdata = 32'd24363;
			41174: outdata = 32'd24362;
			41175: outdata = 32'd24361;
			41176: outdata = 32'd24360;
			41177: outdata = 32'd24359;
			41178: outdata = 32'd24358;
			41179: outdata = 32'd24357;
			41180: outdata = 32'd24356;
			41181: outdata = 32'd24355;
			41182: outdata = 32'd24354;
			41183: outdata = 32'd24353;
			41184: outdata = 32'd24352;
			41185: outdata = 32'd24351;
			41186: outdata = 32'd24350;
			41187: outdata = 32'd24349;
			41188: outdata = 32'd24348;
			41189: outdata = 32'd24347;
			41190: outdata = 32'd24346;
			41191: outdata = 32'd24345;
			41192: outdata = 32'd24344;
			41193: outdata = 32'd24343;
			41194: outdata = 32'd24342;
			41195: outdata = 32'd24341;
			41196: outdata = 32'd24340;
			41197: outdata = 32'd24339;
			41198: outdata = 32'd24338;
			41199: outdata = 32'd24337;
			41200: outdata = 32'd24336;
			41201: outdata = 32'd24335;
			41202: outdata = 32'd24334;
			41203: outdata = 32'd24333;
			41204: outdata = 32'd24332;
			41205: outdata = 32'd24331;
			41206: outdata = 32'd24330;
			41207: outdata = 32'd24329;
			41208: outdata = 32'd24328;
			41209: outdata = 32'd24327;
			41210: outdata = 32'd24326;
			41211: outdata = 32'd24325;
			41212: outdata = 32'd24324;
			41213: outdata = 32'd24323;
			41214: outdata = 32'd24322;
			41215: outdata = 32'd24321;
			41216: outdata = 32'd24320;
			41217: outdata = 32'd24319;
			41218: outdata = 32'd24318;
			41219: outdata = 32'd24317;
			41220: outdata = 32'd24316;
			41221: outdata = 32'd24315;
			41222: outdata = 32'd24314;
			41223: outdata = 32'd24313;
			41224: outdata = 32'd24312;
			41225: outdata = 32'd24311;
			41226: outdata = 32'd24310;
			41227: outdata = 32'd24309;
			41228: outdata = 32'd24308;
			41229: outdata = 32'd24307;
			41230: outdata = 32'd24306;
			41231: outdata = 32'd24305;
			41232: outdata = 32'd24304;
			41233: outdata = 32'd24303;
			41234: outdata = 32'd24302;
			41235: outdata = 32'd24301;
			41236: outdata = 32'd24300;
			41237: outdata = 32'd24299;
			41238: outdata = 32'd24298;
			41239: outdata = 32'd24297;
			41240: outdata = 32'd24296;
			41241: outdata = 32'd24295;
			41242: outdata = 32'd24294;
			41243: outdata = 32'd24293;
			41244: outdata = 32'd24292;
			41245: outdata = 32'd24291;
			41246: outdata = 32'd24290;
			41247: outdata = 32'd24289;
			41248: outdata = 32'd24288;
			41249: outdata = 32'd24287;
			41250: outdata = 32'd24286;
			41251: outdata = 32'd24285;
			41252: outdata = 32'd24284;
			41253: outdata = 32'd24283;
			41254: outdata = 32'd24282;
			41255: outdata = 32'd24281;
			41256: outdata = 32'd24280;
			41257: outdata = 32'd24279;
			41258: outdata = 32'd24278;
			41259: outdata = 32'd24277;
			41260: outdata = 32'd24276;
			41261: outdata = 32'd24275;
			41262: outdata = 32'd24274;
			41263: outdata = 32'd24273;
			41264: outdata = 32'd24272;
			41265: outdata = 32'd24271;
			41266: outdata = 32'd24270;
			41267: outdata = 32'd24269;
			41268: outdata = 32'd24268;
			41269: outdata = 32'd24267;
			41270: outdata = 32'd24266;
			41271: outdata = 32'd24265;
			41272: outdata = 32'd24264;
			41273: outdata = 32'd24263;
			41274: outdata = 32'd24262;
			41275: outdata = 32'd24261;
			41276: outdata = 32'd24260;
			41277: outdata = 32'd24259;
			41278: outdata = 32'd24258;
			41279: outdata = 32'd24257;
			41280: outdata = 32'd24256;
			41281: outdata = 32'd24255;
			41282: outdata = 32'd24254;
			41283: outdata = 32'd24253;
			41284: outdata = 32'd24252;
			41285: outdata = 32'd24251;
			41286: outdata = 32'd24250;
			41287: outdata = 32'd24249;
			41288: outdata = 32'd24248;
			41289: outdata = 32'd24247;
			41290: outdata = 32'd24246;
			41291: outdata = 32'd24245;
			41292: outdata = 32'd24244;
			41293: outdata = 32'd24243;
			41294: outdata = 32'd24242;
			41295: outdata = 32'd24241;
			41296: outdata = 32'd24240;
			41297: outdata = 32'd24239;
			41298: outdata = 32'd24238;
			41299: outdata = 32'd24237;
			41300: outdata = 32'd24236;
			41301: outdata = 32'd24235;
			41302: outdata = 32'd24234;
			41303: outdata = 32'd24233;
			41304: outdata = 32'd24232;
			41305: outdata = 32'd24231;
			41306: outdata = 32'd24230;
			41307: outdata = 32'd24229;
			41308: outdata = 32'd24228;
			41309: outdata = 32'd24227;
			41310: outdata = 32'd24226;
			41311: outdata = 32'd24225;
			41312: outdata = 32'd24224;
			41313: outdata = 32'd24223;
			41314: outdata = 32'd24222;
			41315: outdata = 32'd24221;
			41316: outdata = 32'd24220;
			41317: outdata = 32'd24219;
			41318: outdata = 32'd24218;
			41319: outdata = 32'd24217;
			41320: outdata = 32'd24216;
			41321: outdata = 32'd24215;
			41322: outdata = 32'd24214;
			41323: outdata = 32'd24213;
			41324: outdata = 32'd24212;
			41325: outdata = 32'd24211;
			41326: outdata = 32'd24210;
			41327: outdata = 32'd24209;
			41328: outdata = 32'd24208;
			41329: outdata = 32'd24207;
			41330: outdata = 32'd24206;
			41331: outdata = 32'd24205;
			41332: outdata = 32'd24204;
			41333: outdata = 32'd24203;
			41334: outdata = 32'd24202;
			41335: outdata = 32'd24201;
			41336: outdata = 32'd24200;
			41337: outdata = 32'd24199;
			41338: outdata = 32'd24198;
			41339: outdata = 32'd24197;
			41340: outdata = 32'd24196;
			41341: outdata = 32'd24195;
			41342: outdata = 32'd24194;
			41343: outdata = 32'd24193;
			41344: outdata = 32'd24192;
			41345: outdata = 32'd24191;
			41346: outdata = 32'd24190;
			41347: outdata = 32'd24189;
			41348: outdata = 32'd24188;
			41349: outdata = 32'd24187;
			41350: outdata = 32'd24186;
			41351: outdata = 32'd24185;
			41352: outdata = 32'd24184;
			41353: outdata = 32'd24183;
			41354: outdata = 32'd24182;
			41355: outdata = 32'd24181;
			41356: outdata = 32'd24180;
			41357: outdata = 32'd24179;
			41358: outdata = 32'd24178;
			41359: outdata = 32'd24177;
			41360: outdata = 32'd24176;
			41361: outdata = 32'd24175;
			41362: outdata = 32'd24174;
			41363: outdata = 32'd24173;
			41364: outdata = 32'd24172;
			41365: outdata = 32'd24171;
			41366: outdata = 32'd24170;
			41367: outdata = 32'd24169;
			41368: outdata = 32'd24168;
			41369: outdata = 32'd24167;
			41370: outdata = 32'd24166;
			41371: outdata = 32'd24165;
			41372: outdata = 32'd24164;
			41373: outdata = 32'd24163;
			41374: outdata = 32'd24162;
			41375: outdata = 32'd24161;
			41376: outdata = 32'd24160;
			41377: outdata = 32'd24159;
			41378: outdata = 32'd24158;
			41379: outdata = 32'd24157;
			41380: outdata = 32'd24156;
			41381: outdata = 32'd24155;
			41382: outdata = 32'd24154;
			41383: outdata = 32'd24153;
			41384: outdata = 32'd24152;
			41385: outdata = 32'd24151;
			41386: outdata = 32'd24150;
			41387: outdata = 32'd24149;
			41388: outdata = 32'd24148;
			41389: outdata = 32'd24147;
			41390: outdata = 32'd24146;
			41391: outdata = 32'd24145;
			41392: outdata = 32'd24144;
			41393: outdata = 32'd24143;
			41394: outdata = 32'd24142;
			41395: outdata = 32'd24141;
			41396: outdata = 32'd24140;
			41397: outdata = 32'd24139;
			41398: outdata = 32'd24138;
			41399: outdata = 32'd24137;
			41400: outdata = 32'd24136;
			41401: outdata = 32'd24135;
			41402: outdata = 32'd24134;
			41403: outdata = 32'd24133;
			41404: outdata = 32'd24132;
			41405: outdata = 32'd24131;
			41406: outdata = 32'd24130;
			41407: outdata = 32'd24129;
			41408: outdata = 32'd24128;
			41409: outdata = 32'd24127;
			41410: outdata = 32'd24126;
			41411: outdata = 32'd24125;
			41412: outdata = 32'd24124;
			41413: outdata = 32'd24123;
			41414: outdata = 32'd24122;
			41415: outdata = 32'd24121;
			41416: outdata = 32'd24120;
			41417: outdata = 32'd24119;
			41418: outdata = 32'd24118;
			41419: outdata = 32'd24117;
			41420: outdata = 32'd24116;
			41421: outdata = 32'd24115;
			41422: outdata = 32'd24114;
			41423: outdata = 32'd24113;
			41424: outdata = 32'd24112;
			41425: outdata = 32'd24111;
			41426: outdata = 32'd24110;
			41427: outdata = 32'd24109;
			41428: outdata = 32'd24108;
			41429: outdata = 32'd24107;
			41430: outdata = 32'd24106;
			41431: outdata = 32'd24105;
			41432: outdata = 32'd24104;
			41433: outdata = 32'd24103;
			41434: outdata = 32'd24102;
			41435: outdata = 32'd24101;
			41436: outdata = 32'd24100;
			41437: outdata = 32'd24099;
			41438: outdata = 32'd24098;
			41439: outdata = 32'd24097;
			41440: outdata = 32'd24096;
			41441: outdata = 32'd24095;
			41442: outdata = 32'd24094;
			41443: outdata = 32'd24093;
			41444: outdata = 32'd24092;
			41445: outdata = 32'd24091;
			41446: outdata = 32'd24090;
			41447: outdata = 32'd24089;
			41448: outdata = 32'd24088;
			41449: outdata = 32'd24087;
			41450: outdata = 32'd24086;
			41451: outdata = 32'd24085;
			41452: outdata = 32'd24084;
			41453: outdata = 32'd24083;
			41454: outdata = 32'd24082;
			41455: outdata = 32'd24081;
			41456: outdata = 32'd24080;
			41457: outdata = 32'd24079;
			41458: outdata = 32'd24078;
			41459: outdata = 32'd24077;
			41460: outdata = 32'd24076;
			41461: outdata = 32'd24075;
			41462: outdata = 32'd24074;
			41463: outdata = 32'd24073;
			41464: outdata = 32'd24072;
			41465: outdata = 32'd24071;
			41466: outdata = 32'd24070;
			41467: outdata = 32'd24069;
			41468: outdata = 32'd24068;
			41469: outdata = 32'd24067;
			41470: outdata = 32'd24066;
			41471: outdata = 32'd24065;
			41472: outdata = 32'd24064;
			41473: outdata = 32'd24063;
			41474: outdata = 32'd24062;
			41475: outdata = 32'd24061;
			41476: outdata = 32'd24060;
			41477: outdata = 32'd24059;
			41478: outdata = 32'd24058;
			41479: outdata = 32'd24057;
			41480: outdata = 32'd24056;
			41481: outdata = 32'd24055;
			41482: outdata = 32'd24054;
			41483: outdata = 32'd24053;
			41484: outdata = 32'd24052;
			41485: outdata = 32'd24051;
			41486: outdata = 32'd24050;
			41487: outdata = 32'd24049;
			41488: outdata = 32'd24048;
			41489: outdata = 32'd24047;
			41490: outdata = 32'd24046;
			41491: outdata = 32'd24045;
			41492: outdata = 32'd24044;
			41493: outdata = 32'd24043;
			41494: outdata = 32'd24042;
			41495: outdata = 32'd24041;
			41496: outdata = 32'd24040;
			41497: outdata = 32'd24039;
			41498: outdata = 32'd24038;
			41499: outdata = 32'd24037;
			41500: outdata = 32'd24036;
			41501: outdata = 32'd24035;
			41502: outdata = 32'd24034;
			41503: outdata = 32'd24033;
			41504: outdata = 32'd24032;
			41505: outdata = 32'd24031;
			41506: outdata = 32'd24030;
			41507: outdata = 32'd24029;
			41508: outdata = 32'd24028;
			41509: outdata = 32'd24027;
			41510: outdata = 32'd24026;
			41511: outdata = 32'd24025;
			41512: outdata = 32'd24024;
			41513: outdata = 32'd24023;
			41514: outdata = 32'd24022;
			41515: outdata = 32'd24021;
			41516: outdata = 32'd24020;
			41517: outdata = 32'd24019;
			41518: outdata = 32'd24018;
			41519: outdata = 32'd24017;
			41520: outdata = 32'd24016;
			41521: outdata = 32'd24015;
			41522: outdata = 32'd24014;
			41523: outdata = 32'd24013;
			41524: outdata = 32'd24012;
			41525: outdata = 32'd24011;
			41526: outdata = 32'd24010;
			41527: outdata = 32'd24009;
			41528: outdata = 32'd24008;
			41529: outdata = 32'd24007;
			41530: outdata = 32'd24006;
			41531: outdata = 32'd24005;
			41532: outdata = 32'd24004;
			41533: outdata = 32'd24003;
			41534: outdata = 32'd24002;
			41535: outdata = 32'd24001;
			41536: outdata = 32'd24000;
			41537: outdata = 32'd23999;
			41538: outdata = 32'd23998;
			41539: outdata = 32'd23997;
			41540: outdata = 32'd23996;
			41541: outdata = 32'd23995;
			41542: outdata = 32'd23994;
			41543: outdata = 32'd23993;
			41544: outdata = 32'd23992;
			41545: outdata = 32'd23991;
			41546: outdata = 32'd23990;
			41547: outdata = 32'd23989;
			41548: outdata = 32'd23988;
			41549: outdata = 32'd23987;
			41550: outdata = 32'd23986;
			41551: outdata = 32'd23985;
			41552: outdata = 32'd23984;
			41553: outdata = 32'd23983;
			41554: outdata = 32'd23982;
			41555: outdata = 32'd23981;
			41556: outdata = 32'd23980;
			41557: outdata = 32'd23979;
			41558: outdata = 32'd23978;
			41559: outdata = 32'd23977;
			41560: outdata = 32'd23976;
			41561: outdata = 32'd23975;
			41562: outdata = 32'd23974;
			41563: outdata = 32'd23973;
			41564: outdata = 32'd23972;
			41565: outdata = 32'd23971;
			41566: outdata = 32'd23970;
			41567: outdata = 32'd23969;
			41568: outdata = 32'd23968;
			41569: outdata = 32'd23967;
			41570: outdata = 32'd23966;
			41571: outdata = 32'd23965;
			41572: outdata = 32'd23964;
			41573: outdata = 32'd23963;
			41574: outdata = 32'd23962;
			41575: outdata = 32'd23961;
			41576: outdata = 32'd23960;
			41577: outdata = 32'd23959;
			41578: outdata = 32'd23958;
			41579: outdata = 32'd23957;
			41580: outdata = 32'd23956;
			41581: outdata = 32'd23955;
			41582: outdata = 32'd23954;
			41583: outdata = 32'd23953;
			41584: outdata = 32'd23952;
			41585: outdata = 32'd23951;
			41586: outdata = 32'd23950;
			41587: outdata = 32'd23949;
			41588: outdata = 32'd23948;
			41589: outdata = 32'd23947;
			41590: outdata = 32'd23946;
			41591: outdata = 32'd23945;
			41592: outdata = 32'd23944;
			41593: outdata = 32'd23943;
			41594: outdata = 32'd23942;
			41595: outdata = 32'd23941;
			41596: outdata = 32'd23940;
			41597: outdata = 32'd23939;
			41598: outdata = 32'd23938;
			41599: outdata = 32'd23937;
			41600: outdata = 32'd23936;
			41601: outdata = 32'd23935;
			41602: outdata = 32'd23934;
			41603: outdata = 32'd23933;
			41604: outdata = 32'd23932;
			41605: outdata = 32'd23931;
			41606: outdata = 32'd23930;
			41607: outdata = 32'd23929;
			41608: outdata = 32'd23928;
			41609: outdata = 32'd23927;
			41610: outdata = 32'd23926;
			41611: outdata = 32'd23925;
			41612: outdata = 32'd23924;
			41613: outdata = 32'd23923;
			41614: outdata = 32'd23922;
			41615: outdata = 32'd23921;
			41616: outdata = 32'd23920;
			41617: outdata = 32'd23919;
			41618: outdata = 32'd23918;
			41619: outdata = 32'd23917;
			41620: outdata = 32'd23916;
			41621: outdata = 32'd23915;
			41622: outdata = 32'd23914;
			41623: outdata = 32'd23913;
			41624: outdata = 32'd23912;
			41625: outdata = 32'd23911;
			41626: outdata = 32'd23910;
			41627: outdata = 32'd23909;
			41628: outdata = 32'd23908;
			41629: outdata = 32'd23907;
			41630: outdata = 32'd23906;
			41631: outdata = 32'd23905;
			41632: outdata = 32'd23904;
			41633: outdata = 32'd23903;
			41634: outdata = 32'd23902;
			41635: outdata = 32'd23901;
			41636: outdata = 32'd23900;
			41637: outdata = 32'd23899;
			41638: outdata = 32'd23898;
			41639: outdata = 32'd23897;
			41640: outdata = 32'd23896;
			41641: outdata = 32'd23895;
			41642: outdata = 32'd23894;
			41643: outdata = 32'd23893;
			41644: outdata = 32'd23892;
			41645: outdata = 32'd23891;
			41646: outdata = 32'd23890;
			41647: outdata = 32'd23889;
			41648: outdata = 32'd23888;
			41649: outdata = 32'd23887;
			41650: outdata = 32'd23886;
			41651: outdata = 32'd23885;
			41652: outdata = 32'd23884;
			41653: outdata = 32'd23883;
			41654: outdata = 32'd23882;
			41655: outdata = 32'd23881;
			41656: outdata = 32'd23880;
			41657: outdata = 32'd23879;
			41658: outdata = 32'd23878;
			41659: outdata = 32'd23877;
			41660: outdata = 32'd23876;
			41661: outdata = 32'd23875;
			41662: outdata = 32'd23874;
			41663: outdata = 32'd23873;
			41664: outdata = 32'd23872;
			41665: outdata = 32'd23871;
			41666: outdata = 32'd23870;
			41667: outdata = 32'd23869;
			41668: outdata = 32'd23868;
			41669: outdata = 32'd23867;
			41670: outdata = 32'd23866;
			41671: outdata = 32'd23865;
			41672: outdata = 32'd23864;
			41673: outdata = 32'd23863;
			41674: outdata = 32'd23862;
			41675: outdata = 32'd23861;
			41676: outdata = 32'd23860;
			41677: outdata = 32'd23859;
			41678: outdata = 32'd23858;
			41679: outdata = 32'd23857;
			41680: outdata = 32'd23856;
			41681: outdata = 32'd23855;
			41682: outdata = 32'd23854;
			41683: outdata = 32'd23853;
			41684: outdata = 32'd23852;
			41685: outdata = 32'd23851;
			41686: outdata = 32'd23850;
			41687: outdata = 32'd23849;
			41688: outdata = 32'd23848;
			41689: outdata = 32'd23847;
			41690: outdata = 32'd23846;
			41691: outdata = 32'd23845;
			41692: outdata = 32'd23844;
			41693: outdata = 32'd23843;
			41694: outdata = 32'd23842;
			41695: outdata = 32'd23841;
			41696: outdata = 32'd23840;
			41697: outdata = 32'd23839;
			41698: outdata = 32'd23838;
			41699: outdata = 32'd23837;
			41700: outdata = 32'd23836;
			41701: outdata = 32'd23835;
			41702: outdata = 32'd23834;
			41703: outdata = 32'd23833;
			41704: outdata = 32'd23832;
			41705: outdata = 32'd23831;
			41706: outdata = 32'd23830;
			41707: outdata = 32'd23829;
			41708: outdata = 32'd23828;
			41709: outdata = 32'd23827;
			41710: outdata = 32'd23826;
			41711: outdata = 32'd23825;
			41712: outdata = 32'd23824;
			41713: outdata = 32'd23823;
			41714: outdata = 32'd23822;
			41715: outdata = 32'd23821;
			41716: outdata = 32'd23820;
			41717: outdata = 32'd23819;
			41718: outdata = 32'd23818;
			41719: outdata = 32'd23817;
			41720: outdata = 32'd23816;
			41721: outdata = 32'd23815;
			41722: outdata = 32'd23814;
			41723: outdata = 32'd23813;
			41724: outdata = 32'd23812;
			41725: outdata = 32'd23811;
			41726: outdata = 32'd23810;
			41727: outdata = 32'd23809;
			41728: outdata = 32'd23808;
			41729: outdata = 32'd23807;
			41730: outdata = 32'd23806;
			41731: outdata = 32'd23805;
			41732: outdata = 32'd23804;
			41733: outdata = 32'd23803;
			41734: outdata = 32'd23802;
			41735: outdata = 32'd23801;
			41736: outdata = 32'd23800;
			41737: outdata = 32'd23799;
			41738: outdata = 32'd23798;
			41739: outdata = 32'd23797;
			41740: outdata = 32'd23796;
			41741: outdata = 32'd23795;
			41742: outdata = 32'd23794;
			41743: outdata = 32'd23793;
			41744: outdata = 32'd23792;
			41745: outdata = 32'd23791;
			41746: outdata = 32'd23790;
			41747: outdata = 32'd23789;
			41748: outdata = 32'd23788;
			41749: outdata = 32'd23787;
			41750: outdata = 32'd23786;
			41751: outdata = 32'd23785;
			41752: outdata = 32'd23784;
			41753: outdata = 32'd23783;
			41754: outdata = 32'd23782;
			41755: outdata = 32'd23781;
			41756: outdata = 32'd23780;
			41757: outdata = 32'd23779;
			41758: outdata = 32'd23778;
			41759: outdata = 32'd23777;
			41760: outdata = 32'd23776;
			41761: outdata = 32'd23775;
			41762: outdata = 32'd23774;
			41763: outdata = 32'd23773;
			41764: outdata = 32'd23772;
			41765: outdata = 32'd23771;
			41766: outdata = 32'd23770;
			41767: outdata = 32'd23769;
			41768: outdata = 32'd23768;
			41769: outdata = 32'd23767;
			41770: outdata = 32'd23766;
			41771: outdata = 32'd23765;
			41772: outdata = 32'd23764;
			41773: outdata = 32'd23763;
			41774: outdata = 32'd23762;
			41775: outdata = 32'd23761;
			41776: outdata = 32'd23760;
			41777: outdata = 32'd23759;
			41778: outdata = 32'd23758;
			41779: outdata = 32'd23757;
			41780: outdata = 32'd23756;
			41781: outdata = 32'd23755;
			41782: outdata = 32'd23754;
			41783: outdata = 32'd23753;
			41784: outdata = 32'd23752;
			41785: outdata = 32'd23751;
			41786: outdata = 32'd23750;
			41787: outdata = 32'd23749;
			41788: outdata = 32'd23748;
			41789: outdata = 32'd23747;
			41790: outdata = 32'd23746;
			41791: outdata = 32'd23745;
			41792: outdata = 32'd23744;
			41793: outdata = 32'd23743;
			41794: outdata = 32'd23742;
			41795: outdata = 32'd23741;
			41796: outdata = 32'd23740;
			41797: outdata = 32'd23739;
			41798: outdata = 32'd23738;
			41799: outdata = 32'd23737;
			41800: outdata = 32'd23736;
			41801: outdata = 32'd23735;
			41802: outdata = 32'd23734;
			41803: outdata = 32'd23733;
			41804: outdata = 32'd23732;
			41805: outdata = 32'd23731;
			41806: outdata = 32'd23730;
			41807: outdata = 32'd23729;
			41808: outdata = 32'd23728;
			41809: outdata = 32'd23727;
			41810: outdata = 32'd23726;
			41811: outdata = 32'd23725;
			41812: outdata = 32'd23724;
			41813: outdata = 32'd23723;
			41814: outdata = 32'd23722;
			41815: outdata = 32'd23721;
			41816: outdata = 32'd23720;
			41817: outdata = 32'd23719;
			41818: outdata = 32'd23718;
			41819: outdata = 32'd23717;
			41820: outdata = 32'd23716;
			41821: outdata = 32'd23715;
			41822: outdata = 32'd23714;
			41823: outdata = 32'd23713;
			41824: outdata = 32'd23712;
			41825: outdata = 32'd23711;
			41826: outdata = 32'd23710;
			41827: outdata = 32'd23709;
			41828: outdata = 32'd23708;
			41829: outdata = 32'd23707;
			41830: outdata = 32'd23706;
			41831: outdata = 32'd23705;
			41832: outdata = 32'd23704;
			41833: outdata = 32'd23703;
			41834: outdata = 32'd23702;
			41835: outdata = 32'd23701;
			41836: outdata = 32'd23700;
			41837: outdata = 32'd23699;
			41838: outdata = 32'd23698;
			41839: outdata = 32'd23697;
			41840: outdata = 32'd23696;
			41841: outdata = 32'd23695;
			41842: outdata = 32'd23694;
			41843: outdata = 32'd23693;
			41844: outdata = 32'd23692;
			41845: outdata = 32'd23691;
			41846: outdata = 32'd23690;
			41847: outdata = 32'd23689;
			41848: outdata = 32'd23688;
			41849: outdata = 32'd23687;
			41850: outdata = 32'd23686;
			41851: outdata = 32'd23685;
			41852: outdata = 32'd23684;
			41853: outdata = 32'd23683;
			41854: outdata = 32'd23682;
			41855: outdata = 32'd23681;
			41856: outdata = 32'd23680;
			41857: outdata = 32'd23679;
			41858: outdata = 32'd23678;
			41859: outdata = 32'd23677;
			41860: outdata = 32'd23676;
			41861: outdata = 32'd23675;
			41862: outdata = 32'd23674;
			41863: outdata = 32'd23673;
			41864: outdata = 32'd23672;
			41865: outdata = 32'd23671;
			41866: outdata = 32'd23670;
			41867: outdata = 32'd23669;
			41868: outdata = 32'd23668;
			41869: outdata = 32'd23667;
			41870: outdata = 32'd23666;
			41871: outdata = 32'd23665;
			41872: outdata = 32'd23664;
			41873: outdata = 32'd23663;
			41874: outdata = 32'd23662;
			41875: outdata = 32'd23661;
			41876: outdata = 32'd23660;
			41877: outdata = 32'd23659;
			41878: outdata = 32'd23658;
			41879: outdata = 32'd23657;
			41880: outdata = 32'd23656;
			41881: outdata = 32'd23655;
			41882: outdata = 32'd23654;
			41883: outdata = 32'd23653;
			41884: outdata = 32'd23652;
			41885: outdata = 32'd23651;
			41886: outdata = 32'd23650;
			41887: outdata = 32'd23649;
			41888: outdata = 32'd23648;
			41889: outdata = 32'd23647;
			41890: outdata = 32'd23646;
			41891: outdata = 32'd23645;
			41892: outdata = 32'd23644;
			41893: outdata = 32'd23643;
			41894: outdata = 32'd23642;
			41895: outdata = 32'd23641;
			41896: outdata = 32'd23640;
			41897: outdata = 32'd23639;
			41898: outdata = 32'd23638;
			41899: outdata = 32'd23637;
			41900: outdata = 32'd23636;
			41901: outdata = 32'd23635;
			41902: outdata = 32'd23634;
			41903: outdata = 32'd23633;
			41904: outdata = 32'd23632;
			41905: outdata = 32'd23631;
			41906: outdata = 32'd23630;
			41907: outdata = 32'd23629;
			41908: outdata = 32'd23628;
			41909: outdata = 32'd23627;
			41910: outdata = 32'd23626;
			41911: outdata = 32'd23625;
			41912: outdata = 32'd23624;
			41913: outdata = 32'd23623;
			41914: outdata = 32'd23622;
			41915: outdata = 32'd23621;
			41916: outdata = 32'd23620;
			41917: outdata = 32'd23619;
			41918: outdata = 32'd23618;
			41919: outdata = 32'd23617;
			41920: outdata = 32'd23616;
			41921: outdata = 32'd23615;
			41922: outdata = 32'd23614;
			41923: outdata = 32'd23613;
			41924: outdata = 32'd23612;
			41925: outdata = 32'd23611;
			41926: outdata = 32'd23610;
			41927: outdata = 32'd23609;
			41928: outdata = 32'd23608;
			41929: outdata = 32'd23607;
			41930: outdata = 32'd23606;
			41931: outdata = 32'd23605;
			41932: outdata = 32'd23604;
			41933: outdata = 32'd23603;
			41934: outdata = 32'd23602;
			41935: outdata = 32'd23601;
			41936: outdata = 32'd23600;
			41937: outdata = 32'd23599;
			41938: outdata = 32'd23598;
			41939: outdata = 32'd23597;
			41940: outdata = 32'd23596;
			41941: outdata = 32'd23595;
			41942: outdata = 32'd23594;
			41943: outdata = 32'd23593;
			41944: outdata = 32'd23592;
			41945: outdata = 32'd23591;
			41946: outdata = 32'd23590;
			41947: outdata = 32'd23589;
			41948: outdata = 32'd23588;
			41949: outdata = 32'd23587;
			41950: outdata = 32'd23586;
			41951: outdata = 32'd23585;
			41952: outdata = 32'd23584;
			41953: outdata = 32'd23583;
			41954: outdata = 32'd23582;
			41955: outdata = 32'd23581;
			41956: outdata = 32'd23580;
			41957: outdata = 32'd23579;
			41958: outdata = 32'd23578;
			41959: outdata = 32'd23577;
			41960: outdata = 32'd23576;
			41961: outdata = 32'd23575;
			41962: outdata = 32'd23574;
			41963: outdata = 32'd23573;
			41964: outdata = 32'd23572;
			41965: outdata = 32'd23571;
			41966: outdata = 32'd23570;
			41967: outdata = 32'd23569;
			41968: outdata = 32'd23568;
			41969: outdata = 32'd23567;
			41970: outdata = 32'd23566;
			41971: outdata = 32'd23565;
			41972: outdata = 32'd23564;
			41973: outdata = 32'd23563;
			41974: outdata = 32'd23562;
			41975: outdata = 32'd23561;
			41976: outdata = 32'd23560;
			41977: outdata = 32'd23559;
			41978: outdata = 32'd23558;
			41979: outdata = 32'd23557;
			41980: outdata = 32'd23556;
			41981: outdata = 32'd23555;
			41982: outdata = 32'd23554;
			41983: outdata = 32'd23553;
			41984: outdata = 32'd23552;
			41985: outdata = 32'd23551;
			41986: outdata = 32'd23550;
			41987: outdata = 32'd23549;
			41988: outdata = 32'd23548;
			41989: outdata = 32'd23547;
			41990: outdata = 32'd23546;
			41991: outdata = 32'd23545;
			41992: outdata = 32'd23544;
			41993: outdata = 32'd23543;
			41994: outdata = 32'd23542;
			41995: outdata = 32'd23541;
			41996: outdata = 32'd23540;
			41997: outdata = 32'd23539;
			41998: outdata = 32'd23538;
			41999: outdata = 32'd23537;
			42000: outdata = 32'd23536;
			42001: outdata = 32'd23535;
			42002: outdata = 32'd23534;
			42003: outdata = 32'd23533;
			42004: outdata = 32'd23532;
			42005: outdata = 32'd23531;
			42006: outdata = 32'd23530;
			42007: outdata = 32'd23529;
			42008: outdata = 32'd23528;
			42009: outdata = 32'd23527;
			42010: outdata = 32'd23526;
			42011: outdata = 32'd23525;
			42012: outdata = 32'd23524;
			42013: outdata = 32'd23523;
			42014: outdata = 32'd23522;
			42015: outdata = 32'd23521;
			42016: outdata = 32'd23520;
			42017: outdata = 32'd23519;
			42018: outdata = 32'd23518;
			42019: outdata = 32'd23517;
			42020: outdata = 32'd23516;
			42021: outdata = 32'd23515;
			42022: outdata = 32'd23514;
			42023: outdata = 32'd23513;
			42024: outdata = 32'd23512;
			42025: outdata = 32'd23511;
			42026: outdata = 32'd23510;
			42027: outdata = 32'd23509;
			42028: outdata = 32'd23508;
			42029: outdata = 32'd23507;
			42030: outdata = 32'd23506;
			42031: outdata = 32'd23505;
			42032: outdata = 32'd23504;
			42033: outdata = 32'd23503;
			42034: outdata = 32'd23502;
			42035: outdata = 32'd23501;
			42036: outdata = 32'd23500;
			42037: outdata = 32'd23499;
			42038: outdata = 32'd23498;
			42039: outdata = 32'd23497;
			42040: outdata = 32'd23496;
			42041: outdata = 32'd23495;
			42042: outdata = 32'd23494;
			42043: outdata = 32'd23493;
			42044: outdata = 32'd23492;
			42045: outdata = 32'd23491;
			42046: outdata = 32'd23490;
			42047: outdata = 32'd23489;
			42048: outdata = 32'd23488;
			42049: outdata = 32'd23487;
			42050: outdata = 32'd23486;
			42051: outdata = 32'd23485;
			42052: outdata = 32'd23484;
			42053: outdata = 32'd23483;
			42054: outdata = 32'd23482;
			42055: outdata = 32'd23481;
			42056: outdata = 32'd23480;
			42057: outdata = 32'd23479;
			42058: outdata = 32'd23478;
			42059: outdata = 32'd23477;
			42060: outdata = 32'd23476;
			42061: outdata = 32'd23475;
			42062: outdata = 32'd23474;
			42063: outdata = 32'd23473;
			42064: outdata = 32'd23472;
			42065: outdata = 32'd23471;
			42066: outdata = 32'd23470;
			42067: outdata = 32'd23469;
			42068: outdata = 32'd23468;
			42069: outdata = 32'd23467;
			42070: outdata = 32'd23466;
			42071: outdata = 32'd23465;
			42072: outdata = 32'd23464;
			42073: outdata = 32'd23463;
			42074: outdata = 32'd23462;
			42075: outdata = 32'd23461;
			42076: outdata = 32'd23460;
			42077: outdata = 32'd23459;
			42078: outdata = 32'd23458;
			42079: outdata = 32'd23457;
			42080: outdata = 32'd23456;
			42081: outdata = 32'd23455;
			42082: outdata = 32'd23454;
			42083: outdata = 32'd23453;
			42084: outdata = 32'd23452;
			42085: outdata = 32'd23451;
			42086: outdata = 32'd23450;
			42087: outdata = 32'd23449;
			42088: outdata = 32'd23448;
			42089: outdata = 32'd23447;
			42090: outdata = 32'd23446;
			42091: outdata = 32'd23445;
			42092: outdata = 32'd23444;
			42093: outdata = 32'd23443;
			42094: outdata = 32'd23442;
			42095: outdata = 32'd23441;
			42096: outdata = 32'd23440;
			42097: outdata = 32'd23439;
			42098: outdata = 32'd23438;
			42099: outdata = 32'd23437;
			42100: outdata = 32'd23436;
			42101: outdata = 32'd23435;
			42102: outdata = 32'd23434;
			42103: outdata = 32'd23433;
			42104: outdata = 32'd23432;
			42105: outdata = 32'd23431;
			42106: outdata = 32'd23430;
			42107: outdata = 32'd23429;
			42108: outdata = 32'd23428;
			42109: outdata = 32'd23427;
			42110: outdata = 32'd23426;
			42111: outdata = 32'd23425;
			42112: outdata = 32'd23424;
			42113: outdata = 32'd23423;
			42114: outdata = 32'd23422;
			42115: outdata = 32'd23421;
			42116: outdata = 32'd23420;
			42117: outdata = 32'd23419;
			42118: outdata = 32'd23418;
			42119: outdata = 32'd23417;
			42120: outdata = 32'd23416;
			42121: outdata = 32'd23415;
			42122: outdata = 32'd23414;
			42123: outdata = 32'd23413;
			42124: outdata = 32'd23412;
			42125: outdata = 32'd23411;
			42126: outdata = 32'd23410;
			42127: outdata = 32'd23409;
			42128: outdata = 32'd23408;
			42129: outdata = 32'd23407;
			42130: outdata = 32'd23406;
			42131: outdata = 32'd23405;
			42132: outdata = 32'd23404;
			42133: outdata = 32'd23403;
			42134: outdata = 32'd23402;
			42135: outdata = 32'd23401;
			42136: outdata = 32'd23400;
			42137: outdata = 32'd23399;
			42138: outdata = 32'd23398;
			42139: outdata = 32'd23397;
			42140: outdata = 32'd23396;
			42141: outdata = 32'd23395;
			42142: outdata = 32'd23394;
			42143: outdata = 32'd23393;
			42144: outdata = 32'd23392;
			42145: outdata = 32'd23391;
			42146: outdata = 32'd23390;
			42147: outdata = 32'd23389;
			42148: outdata = 32'd23388;
			42149: outdata = 32'd23387;
			42150: outdata = 32'd23386;
			42151: outdata = 32'd23385;
			42152: outdata = 32'd23384;
			42153: outdata = 32'd23383;
			42154: outdata = 32'd23382;
			42155: outdata = 32'd23381;
			42156: outdata = 32'd23380;
			42157: outdata = 32'd23379;
			42158: outdata = 32'd23378;
			42159: outdata = 32'd23377;
			42160: outdata = 32'd23376;
			42161: outdata = 32'd23375;
			42162: outdata = 32'd23374;
			42163: outdata = 32'd23373;
			42164: outdata = 32'd23372;
			42165: outdata = 32'd23371;
			42166: outdata = 32'd23370;
			42167: outdata = 32'd23369;
			42168: outdata = 32'd23368;
			42169: outdata = 32'd23367;
			42170: outdata = 32'd23366;
			42171: outdata = 32'd23365;
			42172: outdata = 32'd23364;
			42173: outdata = 32'd23363;
			42174: outdata = 32'd23362;
			42175: outdata = 32'd23361;
			42176: outdata = 32'd23360;
			42177: outdata = 32'd23359;
			42178: outdata = 32'd23358;
			42179: outdata = 32'd23357;
			42180: outdata = 32'd23356;
			42181: outdata = 32'd23355;
			42182: outdata = 32'd23354;
			42183: outdata = 32'd23353;
			42184: outdata = 32'd23352;
			42185: outdata = 32'd23351;
			42186: outdata = 32'd23350;
			42187: outdata = 32'd23349;
			42188: outdata = 32'd23348;
			42189: outdata = 32'd23347;
			42190: outdata = 32'd23346;
			42191: outdata = 32'd23345;
			42192: outdata = 32'd23344;
			42193: outdata = 32'd23343;
			42194: outdata = 32'd23342;
			42195: outdata = 32'd23341;
			42196: outdata = 32'd23340;
			42197: outdata = 32'd23339;
			42198: outdata = 32'd23338;
			42199: outdata = 32'd23337;
			42200: outdata = 32'd23336;
			42201: outdata = 32'd23335;
			42202: outdata = 32'd23334;
			42203: outdata = 32'd23333;
			42204: outdata = 32'd23332;
			42205: outdata = 32'd23331;
			42206: outdata = 32'd23330;
			42207: outdata = 32'd23329;
			42208: outdata = 32'd23328;
			42209: outdata = 32'd23327;
			42210: outdata = 32'd23326;
			42211: outdata = 32'd23325;
			42212: outdata = 32'd23324;
			42213: outdata = 32'd23323;
			42214: outdata = 32'd23322;
			42215: outdata = 32'd23321;
			42216: outdata = 32'd23320;
			42217: outdata = 32'd23319;
			42218: outdata = 32'd23318;
			42219: outdata = 32'd23317;
			42220: outdata = 32'd23316;
			42221: outdata = 32'd23315;
			42222: outdata = 32'd23314;
			42223: outdata = 32'd23313;
			42224: outdata = 32'd23312;
			42225: outdata = 32'd23311;
			42226: outdata = 32'd23310;
			42227: outdata = 32'd23309;
			42228: outdata = 32'd23308;
			42229: outdata = 32'd23307;
			42230: outdata = 32'd23306;
			42231: outdata = 32'd23305;
			42232: outdata = 32'd23304;
			42233: outdata = 32'd23303;
			42234: outdata = 32'd23302;
			42235: outdata = 32'd23301;
			42236: outdata = 32'd23300;
			42237: outdata = 32'd23299;
			42238: outdata = 32'd23298;
			42239: outdata = 32'd23297;
			42240: outdata = 32'd23296;
			42241: outdata = 32'd23295;
			42242: outdata = 32'd23294;
			42243: outdata = 32'd23293;
			42244: outdata = 32'd23292;
			42245: outdata = 32'd23291;
			42246: outdata = 32'd23290;
			42247: outdata = 32'd23289;
			42248: outdata = 32'd23288;
			42249: outdata = 32'd23287;
			42250: outdata = 32'd23286;
			42251: outdata = 32'd23285;
			42252: outdata = 32'd23284;
			42253: outdata = 32'd23283;
			42254: outdata = 32'd23282;
			42255: outdata = 32'd23281;
			42256: outdata = 32'd23280;
			42257: outdata = 32'd23279;
			42258: outdata = 32'd23278;
			42259: outdata = 32'd23277;
			42260: outdata = 32'd23276;
			42261: outdata = 32'd23275;
			42262: outdata = 32'd23274;
			42263: outdata = 32'd23273;
			42264: outdata = 32'd23272;
			42265: outdata = 32'd23271;
			42266: outdata = 32'd23270;
			42267: outdata = 32'd23269;
			42268: outdata = 32'd23268;
			42269: outdata = 32'd23267;
			42270: outdata = 32'd23266;
			42271: outdata = 32'd23265;
			42272: outdata = 32'd23264;
			42273: outdata = 32'd23263;
			42274: outdata = 32'd23262;
			42275: outdata = 32'd23261;
			42276: outdata = 32'd23260;
			42277: outdata = 32'd23259;
			42278: outdata = 32'd23258;
			42279: outdata = 32'd23257;
			42280: outdata = 32'd23256;
			42281: outdata = 32'd23255;
			42282: outdata = 32'd23254;
			42283: outdata = 32'd23253;
			42284: outdata = 32'd23252;
			42285: outdata = 32'd23251;
			42286: outdata = 32'd23250;
			42287: outdata = 32'd23249;
			42288: outdata = 32'd23248;
			42289: outdata = 32'd23247;
			42290: outdata = 32'd23246;
			42291: outdata = 32'd23245;
			42292: outdata = 32'd23244;
			42293: outdata = 32'd23243;
			42294: outdata = 32'd23242;
			42295: outdata = 32'd23241;
			42296: outdata = 32'd23240;
			42297: outdata = 32'd23239;
			42298: outdata = 32'd23238;
			42299: outdata = 32'd23237;
			42300: outdata = 32'd23236;
			42301: outdata = 32'd23235;
			42302: outdata = 32'd23234;
			42303: outdata = 32'd23233;
			42304: outdata = 32'd23232;
			42305: outdata = 32'd23231;
			42306: outdata = 32'd23230;
			42307: outdata = 32'd23229;
			42308: outdata = 32'd23228;
			42309: outdata = 32'd23227;
			42310: outdata = 32'd23226;
			42311: outdata = 32'd23225;
			42312: outdata = 32'd23224;
			42313: outdata = 32'd23223;
			42314: outdata = 32'd23222;
			42315: outdata = 32'd23221;
			42316: outdata = 32'd23220;
			42317: outdata = 32'd23219;
			42318: outdata = 32'd23218;
			42319: outdata = 32'd23217;
			42320: outdata = 32'd23216;
			42321: outdata = 32'd23215;
			42322: outdata = 32'd23214;
			42323: outdata = 32'd23213;
			42324: outdata = 32'd23212;
			42325: outdata = 32'd23211;
			42326: outdata = 32'd23210;
			42327: outdata = 32'd23209;
			42328: outdata = 32'd23208;
			42329: outdata = 32'd23207;
			42330: outdata = 32'd23206;
			42331: outdata = 32'd23205;
			42332: outdata = 32'd23204;
			42333: outdata = 32'd23203;
			42334: outdata = 32'd23202;
			42335: outdata = 32'd23201;
			42336: outdata = 32'd23200;
			42337: outdata = 32'd23199;
			42338: outdata = 32'd23198;
			42339: outdata = 32'd23197;
			42340: outdata = 32'd23196;
			42341: outdata = 32'd23195;
			42342: outdata = 32'd23194;
			42343: outdata = 32'd23193;
			42344: outdata = 32'd23192;
			42345: outdata = 32'd23191;
			42346: outdata = 32'd23190;
			42347: outdata = 32'd23189;
			42348: outdata = 32'd23188;
			42349: outdata = 32'd23187;
			42350: outdata = 32'd23186;
			42351: outdata = 32'd23185;
			42352: outdata = 32'd23184;
			42353: outdata = 32'd23183;
			42354: outdata = 32'd23182;
			42355: outdata = 32'd23181;
			42356: outdata = 32'd23180;
			42357: outdata = 32'd23179;
			42358: outdata = 32'd23178;
			42359: outdata = 32'd23177;
			42360: outdata = 32'd23176;
			42361: outdata = 32'd23175;
			42362: outdata = 32'd23174;
			42363: outdata = 32'd23173;
			42364: outdata = 32'd23172;
			42365: outdata = 32'd23171;
			42366: outdata = 32'd23170;
			42367: outdata = 32'd23169;
			42368: outdata = 32'd23168;
			42369: outdata = 32'd23167;
			42370: outdata = 32'd23166;
			42371: outdata = 32'd23165;
			42372: outdata = 32'd23164;
			42373: outdata = 32'd23163;
			42374: outdata = 32'd23162;
			42375: outdata = 32'd23161;
			42376: outdata = 32'd23160;
			42377: outdata = 32'd23159;
			42378: outdata = 32'd23158;
			42379: outdata = 32'd23157;
			42380: outdata = 32'd23156;
			42381: outdata = 32'd23155;
			42382: outdata = 32'd23154;
			42383: outdata = 32'd23153;
			42384: outdata = 32'd23152;
			42385: outdata = 32'd23151;
			42386: outdata = 32'd23150;
			42387: outdata = 32'd23149;
			42388: outdata = 32'd23148;
			42389: outdata = 32'd23147;
			42390: outdata = 32'd23146;
			42391: outdata = 32'd23145;
			42392: outdata = 32'd23144;
			42393: outdata = 32'd23143;
			42394: outdata = 32'd23142;
			42395: outdata = 32'd23141;
			42396: outdata = 32'd23140;
			42397: outdata = 32'd23139;
			42398: outdata = 32'd23138;
			42399: outdata = 32'd23137;
			42400: outdata = 32'd23136;
			42401: outdata = 32'd23135;
			42402: outdata = 32'd23134;
			42403: outdata = 32'd23133;
			42404: outdata = 32'd23132;
			42405: outdata = 32'd23131;
			42406: outdata = 32'd23130;
			42407: outdata = 32'd23129;
			42408: outdata = 32'd23128;
			42409: outdata = 32'd23127;
			42410: outdata = 32'd23126;
			42411: outdata = 32'd23125;
			42412: outdata = 32'd23124;
			42413: outdata = 32'd23123;
			42414: outdata = 32'd23122;
			42415: outdata = 32'd23121;
			42416: outdata = 32'd23120;
			42417: outdata = 32'd23119;
			42418: outdata = 32'd23118;
			42419: outdata = 32'd23117;
			42420: outdata = 32'd23116;
			42421: outdata = 32'd23115;
			42422: outdata = 32'd23114;
			42423: outdata = 32'd23113;
			42424: outdata = 32'd23112;
			42425: outdata = 32'd23111;
			42426: outdata = 32'd23110;
			42427: outdata = 32'd23109;
			42428: outdata = 32'd23108;
			42429: outdata = 32'd23107;
			42430: outdata = 32'd23106;
			42431: outdata = 32'd23105;
			42432: outdata = 32'd23104;
			42433: outdata = 32'd23103;
			42434: outdata = 32'd23102;
			42435: outdata = 32'd23101;
			42436: outdata = 32'd23100;
			42437: outdata = 32'd23099;
			42438: outdata = 32'd23098;
			42439: outdata = 32'd23097;
			42440: outdata = 32'd23096;
			42441: outdata = 32'd23095;
			42442: outdata = 32'd23094;
			42443: outdata = 32'd23093;
			42444: outdata = 32'd23092;
			42445: outdata = 32'd23091;
			42446: outdata = 32'd23090;
			42447: outdata = 32'd23089;
			42448: outdata = 32'd23088;
			42449: outdata = 32'd23087;
			42450: outdata = 32'd23086;
			42451: outdata = 32'd23085;
			42452: outdata = 32'd23084;
			42453: outdata = 32'd23083;
			42454: outdata = 32'd23082;
			42455: outdata = 32'd23081;
			42456: outdata = 32'd23080;
			42457: outdata = 32'd23079;
			42458: outdata = 32'd23078;
			42459: outdata = 32'd23077;
			42460: outdata = 32'd23076;
			42461: outdata = 32'd23075;
			42462: outdata = 32'd23074;
			42463: outdata = 32'd23073;
			42464: outdata = 32'd23072;
			42465: outdata = 32'd23071;
			42466: outdata = 32'd23070;
			42467: outdata = 32'd23069;
			42468: outdata = 32'd23068;
			42469: outdata = 32'd23067;
			42470: outdata = 32'd23066;
			42471: outdata = 32'd23065;
			42472: outdata = 32'd23064;
			42473: outdata = 32'd23063;
			42474: outdata = 32'd23062;
			42475: outdata = 32'd23061;
			42476: outdata = 32'd23060;
			42477: outdata = 32'd23059;
			42478: outdata = 32'd23058;
			42479: outdata = 32'd23057;
			42480: outdata = 32'd23056;
			42481: outdata = 32'd23055;
			42482: outdata = 32'd23054;
			42483: outdata = 32'd23053;
			42484: outdata = 32'd23052;
			42485: outdata = 32'd23051;
			42486: outdata = 32'd23050;
			42487: outdata = 32'd23049;
			42488: outdata = 32'd23048;
			42489: outdata = 32'd23047;
			42490: outdata = 32'd23046;
			42491: outdata = 32'd23045;
			42492: outdata = 32'd23044;
			42493: outdata = 32'd23043;
			42494: outdata = 32'd23042;
			42495: outdata = 32'd23041;
			42496: outdata = 32'd23040;
			42497: outdata = 32'd23039;
			42498: outdata = 32'd23038;
			42499: outdata = 32'd23037;
			42500: outdata = 32'd23036;
			42501: outdata = 32'd23035;
			42502: outdata = 32'd23034;
			42503: outdata = 32'd23033;
			42504: outdata = 32'd23032;
			42505: outdata = 32'd23031;
			42506: outdata = 32'd23030;
			42507: outdata = 32'd23029;
			42508: outdata = 32'd23028;
			42509: outdata = 32'd23027;
			42510: outdata = 32'd23026;
			42511: outdata = 32'd23025;
			42512: outdata = 32'd23024;
			42513: outdata = 32'd23023;
			42514: outdata = 32'd23022;
			42515: outdata = 32'd23021;
			42516: outdata = 32'd23020;
			42517: outdata = 32'd23019;
			42518: outdata = 32'd23018;
			42519: outdata = 32'd23017;
			42520: outdata = 32'd23016;
			42521: outdata = 32'd23015;
			42522: outdata = 32'd23014;
			42523: outdata = 32'd23013;
			42524: outdata = 32'd23012;
			42525: outdata = 32'd23011;
			42526: outdata = 32'd23010;
			42527: outdata = 32'd23009;
			42528: outdata = 32'd23008;
			42529: outdata = 32'd23007;
			42530: outdata = 32'd23006;
			42531: outdata = 32'd23005;
			42532: outdata = 32'd23004;
			42533: outdata = 32'd23003;
			42534: outdata = 32'd23002;
			42535: outdata = 32'd23001;
			42536: outdata = 32'd23000;
			42537: outdata = 32'd22999;
			42538: outdata = 32'd22998;
			42539: outdata = 32'd22997;
			42540: outdata = 32'd22996;
			42541: outdata = 32'd22995;
			42542: outdata = 32'd22994;
			42543: outdata = 32'd22993;
			42544: outdata = 32'd22992;
			42545: outdata = 32'd22991;
			42546: outdata = 32'd22990;
			42547: outdata = 32'd22989;
			42548: outdata = 32'd22988;
			42549: outdata = 32'd22987;
			42550: outdata = 32'd22986;
			42551: outdata = 32'd22985;
			42552: outdata = 32'd22984;
			42553: outdata = 32'd22983;
			42554: outdata = 32'd22982;
			42555: outdata = 32'd22981;
			42556: outdata = 32'd22980;
			42557: outdata = 32'd22979;
			42558: outdata = 32'd22978;
			42559: outdata = 32'd22977;
			42560: outdata = 32'd22976;
			42561: outdata = 32'd22975;
			42562: outdata = 32'd22974;
			42563: outdata = 32'd22973;
			42564: outdata = 32'd22972;
			42565: outdata = 32'd22971;
			42566: outdata = 32'd22970;
			42567: outdata = 32'd22969;
			42568: outdata = 32'd22968;
			42569: outdata = 32'd22967;
			42570: outdata = 32'd22966;
			42571: outdata = 32'd22965;
			42572: outdata = 32'd22964;
			42573: outdata = 32'd22963;
			42574: outdata = 32'd22962;
			42575: outdata = 32'd22961;
			42576: outdata = 32'd22960;
			42577: outdata = 32'd22959;
			42578: outdata = 32'd22958;
			42579: outdata = 32'd22957;
			42580: outdata = 32'd22956;
			42581: outdata = 32'd22955;
			42582: outdata = 32'd22954;
			42583: outdata = 32'd22953;
			42584: outdata = 32'd22952;
			42585: outdata = 32'd22951;
			42586: outdata = 32'd22950;
			42587: outdata = 32'd22949;
			42588: outdata = 32'd22948;
			42589: outdata = 32'd22947;
			42590: outdata = 32'd22946;
			42591: outdata = 32'd22945;
			42592: outdata = 32'd22944;
			42593: outdata = 32'd22943;
			42594: outdata = 32'd22942;
			42595: outdata = 32'd22941;
			42596: outdata = 32'd22940;
			42597: outdata = 32'd22939;
			42598: outdata = 32'd22938;
			42599: outdata = 32'd22937;
			42600: outdata = 32'd22936;
			42601: outdata = 32'd22935;
			42602: outdata = 32'd22934;
			42603: outdata = 32'd22933;
			42604: outdata = 32'd22932;
			42605: outdata = 32'd22931;
			42606: outdata = 32'd22930;
			42607: outdata = 32'd22929;
			42608: outdata = 32'd22928;
			42609: outdata = 32'd22927;
			42610: outdata = 32'd22926;
			42611: outdata = 32'd22925;
			42612: outdata = 32'd22924;
			42613: outdata = 32'd22923;
			42614: outdata = 32'd22922;
			42615: outdata = 32'd22921;
			42616: outdata = 32'd22920;
			42617: outdata = 32'd22919;
			42618: outdata = 32'd22918;
			42619: outdata = 32'd22917;
			42620: outdata = 32'd22916;
			42621: outdata = 32'd22915;
			42622: outdata = 32'd22914;
			42623: outdata = 32'd22913;
			42624: outdata = 32'd22912;
			42625: outdata = 32'd22911;
			42626: outdata = 32'd22910;
			42627: outdata = 32'd22909;
			42628: outdata = 32'd22908;
			42629: outdata = 32'd22907;
			42630: outdata = 32'd22906;
			42631: outdata = 32'd22905;
			42632: outdata = 32'd22904;
			42633: outdata = 32'd22903;
			42634: outdata = 32'd22902;
			42635: outdata = 32'd22901;
			42636: outdata = 32'd22900;
			42637: outdata = 32'd22899;
			42638: outdata = 32'd22898;
			42639: outdata = 32'd22897;
			42640: outdata = 32'd22896;
			42641: outdata = 32'd22895;
			42642: outdata = 32'd22894;
			42643: outdata = 32'd22893;
			42644: outdata = 32'd22892;
			42645: outdata = 32'd22891;
			42646: outdata = 32'd22890;
			42647: outdata = 32'd22889;
			42648: outdata = 32'd22888;
			42649: outdata = 32'd22887;
			42650: outdata = 32'd22886;
			42651: outdata = 32'd22885;
			42652: outdata = 32'd22884;
			42653: outdata = 32'd22883;
			42654: outdata = 32'd22882;
			42655: outdata = 32'd22881;
			42656: outdata = 32'd22880;
			42657: outdata = 32'd22879;
			42658: outdata = 32'd22878;
			42659: outdata = 32'd22877;
			42660: outdata = 32'd22876;
			42661: outdata = 32'd22875;
			42662: outdata = 32'd22874;
			42663: outdata = 32'd22873;
			42664: outdata = 32'd22872;
			42665: outdata = 32'd22871;
			42666: outdata = 32'd22870;
			42667: outdata = 32'd22869;
			42668: outdata = 32'd22868;
			42669: outdata = 32'd22867;
			42670: outdata = 32'd22866;
			42671: outdata = 32'd22865;
			42672: outdata = 32'd22864;
			42673: outdata = 32'd22863;
			42674: outdata = 32'd22862;
			42675: outdata = 32'd22861;
			42676: outdata = 32'd22860;
			42677: outdata = 32'd22859;
			42678: outdata = 32'd22858;
			42679: outdata = 32'd22857;
			42680: outdata = 32'd22856;
			42681: outdata = 32'd22855;
			42682: outdata = 32'd22854;
			42683: outdata = 32'd22853;
			42684: outdata = 32'd22852;
			42685: outdata = 32'd22851;
			42686: outdata = 32'd22850;
			42687: outdata = 32'd22849;
			42688: outdata = 32'd22848;
			42689: outdata = 32'd22847;
			42690: outdata = 32'd22846;
			42691: outdata = 32'd22845;
			42692: outdata = 32'd22844;
			42693: outdata = 32'd22843;
			42694: outdata = 32'd22842;
			42695: outdata = 32'd22841;
			42696: outdata = 32'd22840;
			42697: outdata = 32'd22839;
			42698: outdata = 32'd22838;
			42699: outdata = 32'd22837;
			42700: outdata = 32'd22836;
			42701: outdata = 32'd22835;
			42702: outdata = 32'd22834;
			42703: outdata = 32'd22833;
			42704: outdata = 32'd22832;
			42705: outdata = 32'd22831;
			42706: outdata = 32'd22830;
			42707: outdata = 32'd22829;
			42708: outdata = 32'd22828;
			42709: outdata = 32'd22827;
			42710: outdata = 32'd22826;
			42711: outdata = 32'd22825;
			42712: outdata = 32'd22824;
			42713: outdata = 32'd22823;
			42714: outdata = 32'd22822;
			42715: outdata = 32'd22821;
			42716: outdata = 32'd22820;
			42717: outdata = 32'd22819;
			42718: outdata = 32'd22818;
			42719: outdata = 32'd22817;
			42720: outdata = 32'd22816;
			42721: outdata = 32'd22815;
			42722: outdata = 32'd22814;
			42723: outdata = 32'd22813;
			42724: outdata = 32'd22812;
			42725: outdata = 32'd22811;
			42726: outdata = 32'd22810;
			42727: outdata = 32'd22809;
			42728: outdata = 32'd22808;
			42729: outdata = 32'd22807;
			42730: outdata = 32'd22806;
			42731: outdata = 32'd22805;
			42732: outdata = 32'd22804;
			42733: outdata = 32'd22803;
			42734: outdata = 32'd22802;
			42735: outdata = 32'd22801;
			42736: outdata = 32'd22800;
			42737: outdata = 32'd22799;
			42738: outdata = 32'd22798;
			42739: outdata = 32'd22797;
			42740: outdata = 32'd22796;
			42741: outdata = 32'd22795;
			42742: outdata = 32'd22794;
			42743: outdata = 32'd22793;
			42744: outdata = 32'd22792;
			42745: outdata = 32'd22791;
			42746: outdata = 32'd22790;
			42747: outdata = 32'd22789;
			42748: outdata = 32'd22788;
			42749: outdata = 32'd22787;
			42750: outdata = 32'd22786;
			42751: outdata = 32'd22785;
			42752: outdata = 32'd22784;
			42753: outdata = 32'd22783;
			42754: outdata = 32'd22782;
			42755: outdata = 32'd22781;
			42756: outdata = 32'd22780;
			42757: outdata = 32'd22779;
			42758: outdata = 32'd22778;
			42759: outdata = 32'd22777;
			42760: outdata = 32'd22776;
			42761: outdata = 32'd22775;
			42762: outdata = 32'd22774;
			42763: outdata = 32'd22773;
			42764: outdata = 32'd22772;
			42765: outdata = 32'd22771;
			42766: outdata = 32'd22770;
			42767: outdata = 32'd22769;
			42768: outdata = 32'd22768;
			42769: outdata = 32'd22767;
			42770: outdata = 32'd22766;
			42771: outdata = 32'd22765;
			42772: outdata = 32'd22764;
			42773: outdata = 32'd22763;
			42774: outdata = 32'd22762;
			42775: outdata = 32'd22761;
			42776: outdata = 32'd22760;
			42777: outdata = 32'd22759;
			42778: outdata = 32'd22758;
			42779: outdata = 32'd22757;
			42780: outdata = 32'd22756;
			42781: outdata = 32'd22755;
			42782: outdata = 32'd22754;
			42783: outdata = 32'd22753;
			42784: outdata = 32'd22752;
			42785: outdata = 32'd22751;
			42786: outdata = 32'd22750;
			42787: outdata = 32'd22749;
			42788: outdata = 32'd22748;
			42789: outdata = 32'd22747;
			42790: outdata = 32'd22746;
			42791: outdata = 32'd22745;
			42792: outdata = 32'd22744;
			42793: outdata = 32'd22743;
			42794: outdata = 32'd22742;
			42795: outdata = 32'd22741;
			42796: outdata = 32'd22740;
			42797: outdata = 32'd22739;
			42798: outdata = 32'd22738;
			42799: outdata = 32'd22737;
			42800: outdata = 32'd22736;
			42801: outdata = 32'd22735;
			42802: outdata = 32'd22734;
			42803: outdata = 32'd22733;
			42804: outdata = 32'd22732;
			42805: outdata = 32'd22731;
			42806: outdata = 32'd22730;
			42807: outdata = 32'd22729;
			42808: outdata = 32'd22728;
			42809: outdata = 32'd22727;
			42810: outdata = 32'd22726;
			42811: outdata = 32'd22725;
			42812: outdata = 32'd22724;
			42813: outdata = 32'd22723;
			42814: outdata = 32'd22722;
			42815: outdata = 32'd22721;
			42816: outdata = 32'd22720;
			42817: outdata = 32'd22719;
			42818: outdata = 32'd22718;
			42819: outdata = 32'd22717;
			42820: outdata = 32'd22716;
			42821: outdata = 32'd22715;
			42822: outdata = 32'd22714;
			42823: outdata = 32'd22713;
			42824: outdata = 32'd22712;
			42825: outdata = 32'd22711;
			42826: outdata = 32'd22710;
			42827: outdata = 32'd22709;
			42828: outdata = 32'd22708;
			42829: outdata = 32'd22707;
			42830: outdata = 32'd22706;
			42831: outdata = 32'd22705;
			42832: outdata = 32'd22704;
			42833: outdata = 32'd22703;
			42834: outdata = 32'd22702;
			42835: outdata = 32'd22701;
			42836: outdata = 32'd22700;
			42837: outdata = 32'd22699;
			42838: outdata = 32'd22698;
			42839: outdata = 32'd22697;
			42840: outdata = 32'd22696;
			42841: outdata = 32'd22695;
			42842: outdata = 32'd22694;
			42843: outdata = 32'd22693;
			42844: outdata = 32'd22692;
			42845: outdata = 32'd22691;
			42846: outdata = 32'd22690;
			42847: outdata = 32'd22689;
			42848: outdata = 32'd22688;
			42849: outdata = 32'd22687;
			42850: outdata = 32'd22686;
			42851: outdata = 32'd22685;
			42852: outdata = 32'd22684;
			42853: outdata = 32'd22683;
			42854: outdata = 32'd22682;
			42855: outdata = 32'd22681;
			42856: outdata = 32'd22680;
			42857: outdata = 32'd22679;
			42858: outdata = 32'd22678;
			42859: outdata = 32'd22677;
			42860: outdata = 32'd22676;
			42861: outdata = 32'd22675;
			42862: outdata = 32'd22674;
			42863: outdata = 32'd22673;
			42864: outdata = 32'd22672;
			42865: outdata = 32'd22671;
			42866: outdata = 32'd22670;
			42867: outdata = 32'd22669;
			42868: outdata = 32'd22668;
			42869: outdata = 32'd22667;
			42870: outdata = 32'd22666;
			42871: outdata = 32'd22665;
			42872: outdata = 32'd22664;
			42873: outdata = 32'd22663;
			42874: outdata = 32'd22662;
			42875: outdata = 32'd22661;
			42876: outdata = 32'd22660;
			42877: outdata = 32'd22659;
			42878: outdata = 32'd22658;
			42879: outdata = 32'd22657;
			42880: outdata = 32'd22656;
			42881: outdata = 32'd22655;
			42882: outdata = 32'd22654;
			42883: outdata = 32'd22653;
			42884: outdata = 32'd22652;
			42885: outdata = 32'd22651;
			42886: outdata = 32'd22650;
			42887: outdata = 32'd22649;
			42888: outdata = 32'd22648;
			42889: outdata = 32'd22647;
			42890: outdata = 32'd22646;
			42891: outdata = 32'd22645;
			42892: outdata = 32'd22644;
			42893: outdata = 32'd22643;
			42894: outdata = 32'd22642;
			42895: outdata = 32'd22641;
			42896: outdata = 32'd22640;
			42897: outdata = 32'd22639;
			42898: outdata = 32'd22638;
			42899: outdata = 32'd22637;
			42900: outdata = 32'd22636;
			42901: outdata = 32'd22635;
			42902: outdata = 32'd22634;
			42903: outdata = 32'd22633;
			42904: outdata = 32'd22632;
			42905: outdata = 32'd22631;
			42906: outdata = 32'd22630;
			42907: outdata = 32'd22629;
			42908: outdata = 32'd22628;
			42909: outdata = 32'd22627;
			42910: outdata = 32'd22626;
			42911: outdata = 32'd22625;
			42912: outdata = 32'd22624;
			42913: outdata = 32'd22623;
			42914: outdata = 32'd22622;
			42915: outdata = 32'd22621;
			42916: outdata = 32'd22620;
			42917: outdata = 32'd22619;
			42918: outdata = 32'd22618;
			42919: outdata = 32'd22617;
			42920: outdata = 32'd22616;
			42921: outdata = 32'd22615;
			42922: outdata = 32'd22614;
			42923: outdata = 32'd22613;
			42924: outdata = 32'd22612;
			42925: outdata = 32'd22611;
			42926: outdata = 32'd22610;
			42927: outdata = 32'd22609;
			42928: outdata = 32'd22608;
			42929: outdata = 32'd22607;
			42930: outdata = 32'd22606;
			42931: outdata = 32'd22605;
			42932: outdata = 32'd22604;
			42933: outdata = 32'd22603;
			42934: outdata = 32'd22602;
			42935: outdata = 32'd22601;
			42936: outdata = 32'd22600;
			42937: outdata = 32'd22599;
			42938: outdata = 32'd22598;
			42939: outdata = 32'd22597;
			42940: outdata = 32'd22596;
			42941: outdata = 32'd22595;
			42942: outdata = 32'd22594;
			42943: outdata = 32'd22593;
			42944: outdata = 32'd22592;
			42945: outdata = 32'd22591;
			42946: outdata = 32'd22590;
			42947: outdata = 32'd22589;
			42948: outdata = 32'd22588;
			42949: outdata = 32'd22587;
			42950: outdata = 32'd22586;
			42951: outdata = 32'd22585;
			42952: outdata = 32'd22584;
			42953: outdata = 32'd22583;
			42954: outdata = 32'd22582;
			42955: outdata = 32'd22581;
			42956: outdata = 32'd22580;
			42957: outdata = 32'd22579;
			42958: outdata = 32'd22578;
			42959: outdata = 32'd22577;
			42960: outdata = 32'd22576;
			42961: outdata = 32'd22575;
			42962: outdata = 32'd22574;
			42963: outdata = 32'd22573;
			42964: outdata = 32'd22572;
			42965: outdata = 32'd22571;
			42966: outdata = 32'd22570;
			42967: outdata = 32'd22569;
			42968: outdata = 32'd22568;
			42969: outdata = 32'd22567;
			42970: outdata = 32'd22566;
			42971: outdata = 32'd22565;
			42972: outdata = 32'd22564;
			42973: outdata = 32'd22563;
			42974: outdata = 32'd22562;
			42975: outdata = 32'd22561;
			42976: outdata = 32'd22560;
			42977: outdata = 32'd22559;
			42978: outdata = 32'd22558;
			42979: outdata = 32'd22557;
			42980: outdata = 32'd22556;
			42981: outdata = 32'd22555;
			42982: outdata = 32'd22554;
			42983: outdata = 32'd22553;
			42984: outdata = 32'd22552;
			42985: outdata = 32'd22551;
			42986: outdata = 32'd22550;
			42987: outdata = 32'd22549;
			42988: outdata = 32'd22548;
			42989: outdata = 32'd22547;
			42990: outdata = 32'd22546;
			42991: outdata = 32'd22545;
			42992: outdata = 32'd22544;
			42993: outdata = 32'd22543;
			42994: outdata = 32'd22542;
			42995: outdata = 32'd22541;
			42996: outdata = 32'd22540;
			42997: outdata = 32'd22539;
			42998: outdata = 32'd22538;
			42999: outdata = 32'd22537;
			43000: outdata = 32'd22536;
			43001: outdata = 32'd22535;
			43002: outdata = 32'd22534;
			43003: outdata = 32'd22533;
			43004: outdata = 32'd22532;
			43005: outdata = 32'd22531;
			43006: outdata = 32'd22530;
			43007: outdata = 32'd22529;
			43008: outdata = 32'd22528;
			43009: outdata = 32'd22527;
			43010: outdata = 32'd22526;
			43011: outdata = 32'd22525;
			43012: outdata = 32'd22524;
			43013: outdata = 32'd22523;
			43014: outdata = 32'd22522;
			43015: outdata = 32'd22521;
			43016: outdata = 32'd22520;
			43017: outdata = 32'd22519;
			43018: outdata = 32'd22518;
			43019: outdata = 32'd22517;
			43020: outdata = 32'd22516;
			43021: outdata = 32'd22515;
			43022: outdata = 32'd22514;
			43023: outdata = 32'd22513;
			43024: outdata = 32'd22512;
			43025: outdata = 32'd22511;
			43026: outdata = 32'd22510;
			43027: outdata = 32'd22509;
			43028: outdata = 32'd22508;
			43029: outdata = 32'd22507;
			43030: outdata = 32'd22506;
			43031: outdata = 32'd22505;
			43032: outdata = 32'd22504;
			43033: outdata = 32'd22503;
			43034: outdata = 32'd22502;
			43035: outdata = 32'd22501;
			43036: outdata = 32'd22500;
			43037: outdata = 32'd22499;
			43038: outdata = 32'd22498;
			43039: outdata = 32'd22497;
			43040: outdata = 32'd22496;
			43041: outdata = 32'd22495;
			43042: outdata = 32'd22494;
			43043: outdata = 32'd22493;
			43044: outdata = 32'd22492;
			43045: outdata = 32'd22491;
			43046: outdata = 32'd22490;
			43047: outdata = 32'd22489;
			43048: outdata = 32'd22488;
			43049: outdata = 32'd22487;
			43050: outdata = 32'd22486;
			43051: outdata = 32'd22485;
			43052: outdata = 32'd22484;
			43053: outdata = 32'd22483;
			43054: outdata = 32'd22482;
			43055: outdata = 32'd22481;
			43056: outdata = 32'd22480;
			43057: outdata = 32'd22479;
			43058: outdata = 32'd22478;
			43059: outdata = 32'd22477;
			43060: outdata = 32'd22476;
			43061: outdata = 32'd22475;
			43062: outdata = 32'd22474;
			43063: outdata = 32'd22473;
			43064: outdata = 32'd22472;
			43065: outdata = 32'd22471;
			43066: outdata = 32'd22470;
			43067: outdata = 32'd22469;
			43068: outdata = 32'd22468;
			43069: outdata = 32'd22467;
			43070: outdata = 32'd22466;
			43071: outdata = 32'd22465;
			43072: outdata = 32'd22464;
			43073: outdata = 32'd22463;
			43074: outdata = 32'd22462;
			43075: outdata = 32'd22461;
			43076: outdata = 32'd22460;
			43077: outdata = 32'd22459;
			43078: outdata = 32'd22458;
			43079: outdata = 32'd22457;
			43080: outdata = 32'd22456;
			43081: outdata = 32'd22455;
			43082: outdata = 32'd22454;
			43083: outdata = 32'd22453;
			43084: outdata = 32'd22452;
			43085: outdata = 32'd22451;
			43086: outdata = 32'd22450;
			43087: outdata = 32'd22449;
			43088: outdata = 32'd22448;
			43089: outdata = 32'd22447;
			43090: outdata = 32'd22446;
			43091: outdata = 32'd22445;
			43092: outdata = 32'd22444;
			43093: outdata = 32'd22443;
			43094: outdata = 32'd22442;
			43095: outdata = 32'd22441;
			43096: outdata = 32'd22440;
			43097: outdata = 32'd22439;
			43098: outdata = 32'd22438;
			43099: outdata = 32'd22437;
			43100: outdata = 32'd22436;
			43101: outdata = 32'd22435;
			43102: outdata = 32'd22434;
			43103: outdata = 32'd22433;
			43104: outdata = 32'd22432;
			43105: outdata = 32'd22431;
			43106: outdata = 32'd22430;
			43107: outdata = 32'd22429;
			43108: outdata = 32'd22428;
			43109: outdata = 32'd22427;
			43110: outdata = 32'd22426;
			43111: outdata = 32'd22425;
			43112: outdata = 32'd22424;
			43113: outdata = 32'd22423;
			43114: outdata = 32'd22422;
			43115: outdata = 32'd22421;
			43116: outdata = 32'd22420;
			43117: outdata = 32'd22419;
			43118: outdata = 32'd22418;
			43119: outdata = 32'd22417;
			43120: outdata = 32'd22416;
			43121: outdata = 32'd22415;
			43122: outdata = 32'd22414;
			43123: outdata = 32'd22413;
			43124: outdata = 32'd22412;
			43125: outdata = 32'd22411;
			43126: outdata = 32'd22410;
			43127: outdata = 32'd22409;
			43128: outdata = 32'd22408;
			43129: outdata = 32'd22407;
			43130: outdata = 32'd22406;
			43131: outdata = 32'd22405;
			43132: outdata = 32'd22404;
			43133: outdata = 32'd22403;
			43134: outdata = 32'd22402;
			43135: outdata = 32'd22401;
			43136: outdata = 32'd22400;
			43137: outdata = 32'd22399;
			43138: outdata = 32'd22398;
			43139: outdata = 32'd22397;
			43140: outdata = 32'd22396;
			43141: outdata = 32'd22395;
			43142: outdata = 32'd22394;
			43143: outdata = 32'd22393;
			43144: outdata = 32'd22392;
			43145: outdata = 32'd22391;
			43146: outdata = 32'd22390;
			43147: outdata = 32'd22389;
			43148: outdata = 32'd22388;
			43149: outdata = 32'd22387;
			43150: outdata = 32'd22386;
			43151: outdata = 32'd22385;
			43152: outdata = 32'd22384;
			43153: outdata = 32'd22383;
			43154: outdata = 32'd22382;
			43155: outdata = 32'd22381;
			43156: outdata = 32'd22380;
			43157: outdata = 32'd22379;
			43158: outdata = 32'd22378;
			43159: outdata = 32'd22377;
			43160: outdata = 32'd22376;
			43161: outdata = 32'd22375;
			43162: outdata = 32'd22374;
			43163: outdata = 32'd22373;
			43164: outdata = 32'd22372;
			43165: outdata = 32'd22371;
			43166: outdata = 32'd22370;
			43167: outdata = 32'd22369;
			43168: outdata = 32'd22368;
			43169: outdata = 32'd22367;
			43170: outdata = 32'd22366;
			43171: outdata = 32'd22365;
			43172: outdata = 32'd22364;
			43173: outdata = 32'd22363;
			43174: outdata = 32'd22362;
			43175: outdata = 32'd22361;
			43176: outdata = 32'd22360;
			43177: outdata = 32'd22359;
			43178: outdata = 32'd22358;
			43179: outdata = 32'd22357;
			43180: outdata = 32'd22356;
			43181: outdata = 32'd22355;
			43182: outdata = 32'd22354;
			43183: outdata = 32'd22353;
			43184: outdata = 32'd22352;
			43185: outdata = 32'd22351;
			43186: outdata = 32'd22350;
			43187: outdata = 32'd22349;
			43188: outdata = 32'd22348;
			43189: outdata = 32'd22347;
			43190: outdata = 32'd22346;
			43191: outdata = 32'd22345;
			43192: outdata = 32'd22344;
			43193: outdata = 32'd22343;
			43194: outdata = 32'd22342;
			43195: outdata = 32'd22341;
			43196: outdata = 32'd22340;
			43197: outdata = 32'd22339;
			43198: outdata = 32'd22338;
			43199: outdata = 32'd22337;
			43200: outdata = 32'd22336;
			43201: outdata = 32'd22335;
			43202: outdata = 32'd22334;
			43203: outdata = 32'd22333;
			43204: outdata = 32'd22332;
			43205: outdata = 32'd22331;
			43206: outdata = 32'd22330;
			43207: outdata = 32'd22329;
			43208: outdata = 32'd22328;
			43209: outdata = 32'd22327;
			43210: outdata = 32'd22326;
			43211: outdata = 32'd22325;
			43212: outdata = 32'd22324;
			43213: outdata = 32'd22323;
			43214: outdata = 32'd22322;
			43215: outdata = 32'd22321;
			43216: outdata = 32'd22320;
			43217: outdata = 32'd22319;
			43218: outdata = 32'd22318;
			43219: outdata = 32'd22317;
			43220: outdata = 32'd22316;
			43221: outdata = 32'd22315;
			43222: outdata = 32'd22314;
			43223: outdata = 32'd22313;
			43224: outdata = 32'd22312;
			43225: outdata = 32'd22311;
			43226: outdata = 32'd22310;
			43227: outdata = 32'd22309;
			43228: outdata = 32'd22308;
			43229: outdata = 32'd22307;
			43230: outdata = 32'd22306;
			43231: outdata = 32'd22305;
			43232: outdata = 32'd22304;
			43233: outdata = 32'd22303;
			43234: outdata = 32'd22302;
			43235: outdata = 32'd22301;
			43236: outdata = 32'd22300;
			43237: outdata = 32'd22299;
			43238: outdata = 32'd22298;
			43239: outdata = 32'd22297;
			43240: outdata = 32'd22296;
			43241: outdata = 32'd22295;
			43242: outdata = 32'd22294;
			43243: outdata = 32'd22293;
			43244: outdata = 32'd22292;
			43245: outdata = 32'd22291;
			43246: outdata = 32'd22290;
			43247: outdata = 32'd22289;
			43248: outdata = 32'd22288;
			43249: outdata = 32'd22287;
			43250: outdata = 32'd22286;
			43251: outdata = 32'd22285;
			43252: outdata = 32'd22284;
			43253: outdata = 32'd22283;
			43254: outdata = 32'd22282;
			43255: outdata = 32'd22281;
			43256: outdata = 32'd22280;
			43257: outdata = 32'd22279;
			43258: outdata = 32'd22278;
			43259: outdata = 32'd22277;
			43260: outdata = 32'd22276;
			43261: outdata = 32'd22275;
			43262: outdata = 32'd22274;
			43263: outdata = 32'd22273;
			43264: outdata = 32'd22272;
			43265: outdata = 32'd22271;
			43266: outdata = 32'd22270;
			43267: outdata = 32'd22269;
			43268: outdata = 32'd22268;
			43269: outdata = 32'd22267;
			43270: outdata = 32'd22266;
			43271: outdata = 32'd22265;
			43272: outdata = 32'd22264;
			43273: outdata = 32'd22263;
			43274: outdata = 32'd22262;
			43275: outdata = 32'd22261;
			43276: outdata = 32'd22260;
			43277: outdata = 32'd22259;
			43278: outdata = 32'd22258;
			43279: outdata = 32'd22257;
			43280: outdata = 32'd22256;
			43281: outdata = 32'd22255;
			43282: outdata = 32'd22254;
			43283: outdata = 32'd22253;
			43284: outdata = 32'd22252;
			43285: outdata = 32'd22251;
			43286: outdata = 32'd22250;
			43287: outdata = 32'd22249;
			43288: outdata = 32'd22248;
			43289: outdata = 32'd22247;
			43290: outdata = 32'd22246;
			43291: outdata = 32'd22245;
			43292: outdata = 32'd22244;
			43293: outdata = 32'd22243;
			43294: outdata = 32'd22242;
			43295: outdata = 32'd22241;
			43296: outdata = 32'd22240;
			43297: outdata = 32'd22239;
			43298: outdata = 32'd22238;
			43299: outdata = 32'd22237;
			43300: outdata = 32'd22236;
			43301: outdata = 32'd22235;
			43302: outdata = 32'd22234;
			43303: outdata = 32'd22233;
			43304: outdata = 32'd22232;
			43305: outdata = 32'd22231;
			43306: outdata = 32'd22230;
			43307: outdata = 32'd22229;
			43308: outdata = 32'd22228;
			43309: outdata = 32'd22227;
			43310: outdata = 32'd22226;
			43311: outdata = 32'd22225;
			43312: outdata = 32'd22224;
			43313: outdata = 32'd22223;
			43314: outdata = 32'd22222;
			43315: outdata = 32'd22221;
			43316: outdata = 32'd22220;
			43317: outdata = 32'd22219;
			43318: outdata = 32'd22218;
			43319: outdata = 32'd22217;
			43320: outdata = 32'd22216;
			43321: outdata = 32'd22215;
			43322: outdata = 32'd22214;
			43323: outdata = 32'd22213;
			43324: outdata = 32'd22212;
			43325: outdata = 32'd22211;
			43326: outdata = 32'd22210;
			43327: outdata = 32'd22209;
			43328: outdata = 32'd22208;
			43329: outdata = 32'd22207;
			43330: outdata = 32'd22206;
			43331: outdata = 32'd22205;
			43332: outdata = 32'd22204;
			43333: outdata = 32'd22203;
			43334: outdata = 32'd22202;
			43335: outdata = 32'd22201;
			43336: outdata = 32'd22200;
			43337: outdata = 32'd22199;
			43338: outdata = 32'd22198;
			43339: outdata = 32'd22197;
			43340: outdata = 32'd22196;
			43341: outdata = 32'd22195;
			43342: outdata = 32'd22194;
			43343: outdata = 32'd22193;
			43344: outdata = 32'd22192;
			43345: outdata = 32'd22191;
			43346: outdata = 32'd22190;
			43347: outdata = 32'd22189;
			43348: outdata = 32'd22188;
			43349: outdata = 32'd22187;
			43350: outdata = 32'd22186;
			43351: outdata = 32'd22185;
			43352: outdata = 32'd22184;
			43353: outdata = 32'd22183;
			43354: outdata = 32'd22182;
			43355: outdata = 32'd22181;
			43356: outdata = 32'd22180;
			43357: outdata = 32'd22179;
			43358: outdata = 32'd22178;
			43359: outdata = 32'd22177;
			43360: outdata = 32'd22176;
			43361: outdata = 32'd22175;
			43362: outdata = 32'd22174;
			43363: outdata = 32'd22173;
			43364: outdata = 32'd22172;
			43365: outdata = 32'd22171;
			43366: outdata = 32'd22170;
			43367: outdata = 32'd22169;
			43368: outdata = 32'd22168;
			43369: outdata = 32'd22167;
			43370: outdata = 32'd22166;
			43371: outdata = 32'd22165;
			43372: outdata = 32'd22164;
			43373: outdata = 32'd22163;
			43374: outdata = 32'd22162;
			43375: outdata = 32'd22161;
			43376: outdata = 32'd22160;
			43377: outdata = 32'd22159;
			43378: outdata = 32'd22158;
			43379: outdata = 32'd22157;
			43380: outdata = 32'd22156;
			43381: outdata = 32'd22155;
			43382: outdata = 32'd22154;
			43383: outdata = 32'd22153;
			43384: outdata = 32'd22152;
			43385: outdata = 32'd22151;
			43386: outdata = 32'd22150;
			43387: outdata = 32'd22149;
			43388: outdata = 32'd22148;
			43389: outdata = 32'd22147;
			43390: outdata = 32'd22146;
			43391: outdata = 32'd22145;
			43392: outdata = 32'd22144;
			43393: outdata = 32'd22143;
			43394: outdata = 32'd22142;
			43395: outdata = 32'd22141;
			43396: outdata = 32'd22140;
			43397: outdata = 32'd22139;
			43398: outdata = 32'd22138;
			43399: outdata = 32'd22137;
			43400: outdata = 32'd22136;
			43401: outdata = 32'd22135;
			43402: outdata = 32'd22134;
			43403: outdata = 32'd22133;
			43404: outdata = 32'd22132;
			43405: outdata = 32'd22131;
			43406: outdata = 32'd22130;
			43407: outdata = 32'd22129;
			43408: outdata = 32'd22128;
			43409: outdata = 32'd22127;
			43410: outdata = 32'd22126;
			43411: outdata = 32'd22125;
			43412: outdata = 32'd22124;
			43413: outdata = 32'd22123;
			43414: outdata = 32'd22122;
			43415: outdata = 32'd22121;
			43416: outdata = 32'd22120;
			43417: outdata = 32'd22119;
			43418: outdata = 32'd22118;
			43419: outdata = 32'd22117;
			43420: outdata = 32'd22116;
			43421: outdata = 32'd22115;
			43422: outdata = 32'd22114;
			43423: outdata = 32'd22113;
			43424: outdata = 32'd22112;
			43425: outdata = 32'd22111;
			43426: outdata = 32'd22110;
			43427: outdata = 32'd22109;
			43428: outdata = 32'd22108;
			43429: outdata = 32'd22107;
			43430: outdata = 32'd22106;
			43431: outdata = 32'd22105;
			43432: outdata = 32'd22104;
			43433: outdata = 32'd22103;
			43434: outdata = 32'd22102;
			43435: outdata = 32'd22101;
			43436: outdata = 32'd22100;
			43437: outdata = 32'd22099;
			43438: outdata = 32'd22098;
			43439: outdata = 32'd22097;
			43440: outdata = 32'd22096;
			43441: outdata = 32'd22095;
			43442: outdata = 32'd22094;
			43443: outdata = 32'd22093;
			43444: outdata = 32'd22092;
			43445: outdata = 32'd22091;
			43446: outdata = 32'd22090;
			43447: outdata = 32'd22089;
			43448: outdata = 32'd22088;
			43449: outdata = 32'd22087;
			43450: outdata = 32'd22086;
			43451: outdata = 32'd22085;
			43452: outdata = 32'd22084;
			43453: outdata = 32'd22083;
			43454: outdata = 32'd22082;
			43455: outdata = 32'd22081;
			43456: outdata = 32'd22080;
			43457: outdata = 32'd22079;
			43458: outdata = 32'd22078;
			43459: outdata = 32'd22077;
			43460: outdata = 32'd22076;
			43461: outdata = 32'd22075;
			43462: outdata = 32'd22074;
			43463: outdata = 32'd22073;
			43464: outdata = 32'd22072;
			43465: outdata = 32'd22071;
			43466: outdata = 32'd22070;
			43467: outdata = 32'd22069;
			43468: outdata = 32'd22068;
			43469: outdata = 32'd22067;
			43470: outdata = 32'd22066;
			43471: outdata = 32'd22065;
			43472: outdata = 32'd22064;
			43473: outdata = 32'd22063;
			43474: outdata = 32'd22062;
			43475: outdata = 32'd22061;
			43476: outdata = 32'd22060;
			43477: outdata = 32'd22059;
			43478: outdata = 32'd22058;
			43479: outdata = 32'd22057;
			43480: outdata = 32'd22056;
			43481: outdata = 32'd22055;
			43482: outdata = 32'd22054;
			43483: outdata = 32'd22053;
			43484: outdata = 32'd22052;
			43485: outdata = 32'd22051;
			43486: outdata = 32'd22050;
			43487: outdata = 32'd22049;
			43488: outdata = 32'd22048;
			43489: outdata = 32'd22047;
			43490: outdata = 32'd22046;
			43491: outdata = 32'd22045;
			43492: outdata = 32'd22044;
			43493: outdata = 32'd22043;
			43494: outdata = 32'd22042;
			43495: outdata = 32'd22041;
			43496: outdata = 32'd22040;
			43497: outdata = 32'd22039;
			43498: outdata = 32'd22038;
			43499: outdata = 32'd22037;
			43500: outdata = 32'd22036;
			43501: outdata = 32'd22035;
			43502: outdata = 32'd22034;
			43503: outdata = 32'd22033;
			43504: outdata = 32'd22032;
			43505: outdata = 32'd22031;
			43506: outdata = 32'd22030;
			43507: outdata = 32'd22029;
			43508: outdata = 32'd22028;
			43509: outdata = 32'd22027;
			43510: outdata = 32'd22026;
			43511: outdata = 32'd22025;
			43512: outdata = 32'd22024;
			43513: outdata = 32'd22023;
			43514: outdata = 32'd22022;
			43515: outdata = 32'd22021;
			43516: outdata = 32'd22020;
			43517: outdata = 32'd22019;
			43518: outdata = 32'd22018;
			43519: outdata = 32'd22017;
			43520: outdata = 32'd22016;
			43521: outdata = 32'd22015;
			43522: outdata = 32'd22014;
			43523: outdata = 32'd22013;
			43524: outdata = 32'd22012;
			43525: outdata = 32'd22011;
			43526: outdata = 32'd22010;
			43527: outdata = 32'd22009;
			43528: outdata = 32'd22008;
			43529: outdata = 32'd22007;
			43530: outdata = 32'd22006;
			43531: outdata = 32'd22005;
			43532: outdata = 32'd22004;
			43533: outdata = 32'd22003;
			43534: outdata = 32'd22002;
			43535: outdata = 32'd22001;
			43536: outdata = 32'd22000;
			43537: outdata = 32'd21999;
			43538: outdata = 32'd21998;
			43539: outdata = 32'd21997;
			43540: outdata = 32'd21996;
			43541: outdata = 32'd21995;
			43542: outdata = 32'd21994;
			43543: outdata = 32'd21993;
			43544: outdata = 32'd21992;
			43545: outdata = 32'd21991;
			43546: outdata = 32'd21990;
			43547: outdata = 32'd21989;
			43548: outdata = 32'd21988;
			43549: outdata = 32'd21987;
			43550: outdata = 32'd21986;
			43551: outdata = 32'd21985;
			43552: outdata = 32'd21984;
			43553: outdata = 32'd21983;
			43554: outdata = 32'd21982;
			43555: outdata = 32'd21981;
			43556: outdata = 32'd21980;
			43557: outdata = 32'd21979;
			43558: outdata = 32'd21978;
			43559: outdata = 32'd21977;
			43560: outdata = 32'd21976;
			43561: outdata = 32'd21975;
			43562: outdata = 32'd21974;
			43563: outdata = 32'd21973;
			43564: outdata = 32'd21972;
			43565: outdata = 32'd21971;
			43566: outdata = 32'd21970;
			43567: outdata = 32'd21969;
			43568: outdata = 32'd21968;
			43569: outdata = 32'd21967;
			43570: outdata = 32'd21966;
			43571: outdata = 32'd21965;
			43572: outdata = 32'd21964;
			43573: outdata = 32'd21963;
			43574: outdata = 32'd21962;
			43575: outdata = 32'd21961;
			43576: outdata = 32'd21960;
			43577: outdata = 32'd21959;
			43578: outdata = 32'd21958;
			43579: outdata = 32'd21957;
			43580: outdata = 32'd21956;
			43581: outdata = 32'd21955;
			43582: outdata = 32'd21954;
			43583: outdata = 32'd21953;
			43584: outdata = 32'd21952;
			43585: outdata = 32'd21951;
			43586: outdata = 32'd21950;
			43587: outdata = 32'd21949;
			43588: outdata = 32'd21948;
			43589: outdata = 32'd21947;
			43590: outdata = 32'd21946;
			43591: outdata = 32'd21945;
			43592: outdata = 32'd21944;
			43593: outdata = 32'd21943;
			43594: outdata = 32'd21942;
			43595: outdata = 32'd21941;
			43596: outdata = 32'd21940;
			43597: outdata = 32'd21939;
			43598: outdata = 32'd21938;
			43599: outdata = 32'd21937;
			43600: outdata = 32'd21936;
			43601: outdata = 32'd21935;
			43602: outdata = 32'd21934;
			43603: outdata = 32'd21933;
			43604: outdata = 32'd21932;
			43605: outdata = 32'd21931;
			43606: outdata = 32'd21930;
			43607: outdata = 32'd21929;
			43608: outdata = 32'd21928;
			43609: outdata = 32'd21927;
			43610: outdata = 32'd21926;
			43611: outdata = 32'd21925;
			43612: outdata = 32'd21924;
			43613: outdata = 32'd21923;
			43614: outdata = 32'd21922;
			43615: outdata = 32'd21921;
			43616: outdata = 32'd21920;
			43617: outdata = 32'd21919;
			43618: outdata = 32'd21918;
			43619: outdata = 32'd21917;
			43620: outdata = 32'd21916;
			43621: outdata = 32'd21915;
			43622: outdata = 32'd21914;
			43623: outdata = 32'd21913;
			43624: outdata = 32'd21912;
			43625: outdata = 32'd21911;
			43626: outdata = 32'd21910;
			43627: outdata = 32'd21909;
			43628: outdata = 32'd21908;
			43629: outdata = 32'd21907;
			43630: outdata = 32'd21906;
			43631: outdata = 32'd21905;
			43632: outdata = 32'd21904;
			43633: outdata = 32'd21903;
			43634: outdata = 32'd21902;
			43635: outdata = 32'd21901;
			43636: outdata = 32'd21900;
			43637: outdata = 32'd21899;
			43638: outdata = 32'd21898;
			43639: outdata = 32'd21897;
			43640: outdata = 32'd21896;
			43641: outdata = 32'd21895;
			43642: outdata = 32'd21894;
			43643: outdata = 32'd21893;
			43644: outdata = 32'd21892;
			43645: outdata = 32'd21891;
			43646: outdata = 32'd21890;
			43647: outdata = 32'd21889;
			43648: outdata = 32'd21888;
			43649: outdata = 32'd21887;
			43650: outdata = 32'd21886;
			43651: outdata = 32'd21885;
			43652: outdata = 32'd21884;
			43653: outdata = 32'd21883;
			43654: outdata = 32'd21882;
			43655: outdata = 32'd21881;
			43656: outdata = 32'd21880;
			43657: outdata = 32'd21879;
			43658: outdata = 32'd21878;
			43659: outdata = 32'd21877;
			43660: outdata = 32'd21876;
			43661: outdata = 32'd21875;
			43662: outdata = 32'd21874;
			43663: outdata = 32'd21873;
			43664: outdata = 32'd21872;
			43665: outdata = 32'd21871;
			43666: outdata = 32'd21870;
			43667: outdata = 32'd21869;
			43668: outdata = 32'd21868;
			43669: outdata = 32'd21867;
			43670: outdata = 32'd21866;
			43671: outdata = 32'd21865;
			43672: outdata = 32'd21864;
			43673: outdata = 32'd21863;
			43674: outdata = 32'd21862;
			43675: outdata = 32'd21861;
			43676: outdata = 32'd21860;
			43677: outdata = 32'd21859;
			43678: outdata = 32'd21858;
			43679: outdata = 32'd21857;
			43680: outdata = 32'd21856;
			43681: outdata = 32'd21855;
			43682: outdata = 32'd21854;
			43683: outdata = 32'd21853;
			43684: outdata = 32'd21852;
			43685: outdata = 32'd21851;
			43686: outdata = 32'd21850;
			43687: outdata = 32'd21849;
			43688: outdata = 32'd21848;
			43689: outdata = 32'd21847;
			43690: outdata = 32'd21846;
			43691: outdata = 32'd21845;
			43692: outdata = 32'd21844;
			43693: outdata = 32'd21843;
			43694: outdata = 32'd21842;
			43695: outdata = 32'd21841;
			43696: outdata = 32'd21840;
			43697: outdata = 32'd21839;
			43698: outdata = 32'd21838;
			43699: outdata = 32'd21837;
			43700: outdata = 32'd21836;
			43701: outdata = 32'd21835;
			43702: outdata = 32'd21834;
			43703: outdata = 32'd21833;
			43704: outdata = 32'd21832;
			43705: outdata = 32'd21831;
			43706: outdata = 32'd21830;
			43707: outdata = 32'd21829;
			43708: outdata = 32'd21828;
			43709: outdata = 32'd21827;
			43710: outdata = 32'd21826;
			43711: outdata = 32'd21825;
			43712: outdata = 32'd21824;
			43713: outdata = 32'd21823;
			43714: outdata = 32'd21822;
			43715: outdata = 32'd21821;
			43716: outdata = 32'd21820;
			43717: outdata = 32'd21819;
			43718: outdata = 32'd21818;
			43719: outdata = 32'd21817;
			43720: outdata = 32'd21816;
			43721: outdata = 32'd21815;
			43722: outdata = 32'd21814;
			43723: outdata = 32'd21813;
			43724: outdata = 32'd21812;
			43725: outdata = 32'd21811;
			43726: outdata = 32'd21810;
			43727: outdata = 32'd21809;
			43728: outdata = 32'd21808;
			43729: outdata = 32'd21807;
			43730: outdata = 32'd21806;
			43731: outdata = 32'd21805;
			43732: outdata = 32'd21804;
			43733: outdata = 32'd21803;
			43734: outdata = 32'd21802;
			43735: outdata = 32'd21801;
			43736: outdata = 32'd21800;
			43737: outdata = 32'd21799;
			43738: outdata = 32'd21798;
			43739: outdata = 32'd21797;
			43740: outdata = 32'd21796;
			43741: outdata = 32'd21795;
			43742: outdata = 32'd21794;
			43743: outdata = 32'd21793;
			43744: outdata = 32'd21792;
			43745: outdata = 32'd21791;
			43746: outdata = 32'd21790;
			43747: outdata = 32'd21789;
			43748: outdata = 32'd21788;
			43749: outdata = 32'd21787;
			43750: outdata = 32'd21786;
			43751: outdata = 32'd21785;
			43752: outdata = 32'd21784;
			43753: outdata = 32'd21783;
			43754: outdata = 32'd21782;
			43755: outdata = 32'd21781;
			43756: outdata = 32'd21780;
			43757: outdata = 32'd21779;
			43758: outdata = 32'd21778;
			43759: outdata = 32'd21777;
			43760: outdata = 32'd21776;
			43761: outdata = 32'd21775;
			43762: outdata = 32'd21774;
			43763: outdata = 32'd21773;
			43764: outdata = 32'd21772;
			43765: outdata = 32'd21771;
			43766: outdata = 32'd21770;
			43767: outdata = 32'd21769;
			43768: outdata = 32'd21768;
			43769: outdata = 32'd21767;
			43770: outdata = 32'd21766;
			43771: outdata = 32'd21765;
			43772: outdata = 32'd21764;
			43773: outdata = 32'd21763;
			43774: outdata = 32'd21762;
			43775: outdata = 32'd21761;
			43776: outdata = 32'd21760;
			43777: outdata = 32'd21759;
			43778: outdata = 32'd21758;
			43779: outdata = 32'd21757;
			43780: outdata = 32'd21756;
			43781: outdata = 32'd21755;
			43782: outdata = 32'd21754;
			43783: outdata = 32'd21753;
			43784: outdata = 32'd21752;
			43785: outdata = 32'd21751;
			43786: outdata = 32'd21750;
			43787: outdata = 32'd21749;
			43788: outdata = 32'd21748;
			43789: outdata = 32'd21747;
			43790: outdata = 32'd21746;
			43791: outdata = 32'd21745;
			43792: outdata = 32'd21744;
			43793: outdata = 32'd21743;
			43794: outdata = 32'd21742;
			43795: outdata = 32'd21741;
			43796: outdata = 32'd21740;
			43797: outdata = 32'd21739;
			43798: outdata = 32'd21738;
			43799: outdata = 32'd21737;
			43800: outdata = 32'd21736;
			43801: outdata = 32'd21735;
			43802: outdata = 32'd21734;
			43803: outdata = 32'd21733;
			43804: outdata = 32'd21732;
			43805: outdata = 32'd21731;
			43806: outdata = 32'd21730;
			43807: outdata = 32'd21729;
			43808: outdata = 32'd21728;
			43809: outdata = 32'd21727;
			43810: outdata = 32'd21726;
			43811: outdata = 32'd21725;
			43812: outdata = 32'd21724;
			43813: outdata = 32'd21723;
			43814: outdata = 32'd21722;
			43815: outdata = 32'd21721;
			43816: outdata = 32'd21720;
			43817: outdata = 32'd21719;
			43818: outdata = 32'd21718;
			43819: outdata = 32'd21717;
			43820: outdata = 32'd21716;
			43821: outdata = 32'd21715;
			43822: outdata = 32'd21714;
			43823: outdata = 32'd21713;
			43824: outdata = 32'd21712;
			43825: outdata = 32'd21711;
			43826: outdata = 32'd21710;
			43827: outdata = 32'd21709;
			43828: outdata = 32'd21708;
			43829: outdata = 32'd21707;
			43830: outdata = 32'd21706;
			43831: outdata = 32'd21705;
			43832: outdata = 32'd21704;
			43833: outdata = 32'd21703;
			43834: outdata = 32'd21702;
			43835: outdata = 32'd21701;
			43836: outdata = 32'd21700;
			43837: outdata = 32'd21699;
			43838: outdata = 32'd21698;
			43839: outdata = 32'd21697;
			43840: outdata = 32'd21696;
			43841: outdata = 32'd21695;
			43842: outdata = 32'd21694;
			43843: outdata = 32'd21693;
			43844: outdata = 32'd21692;
			43845: outdata = 32'd21691;
			43846: outdata = 32'd21690;
			43847: outdata = 32'd21689;
			43848: outdata = 32'd21688;
			43849: outdata = 32'd21687;
			43850: outdata = 32'd21686;
			43851: outdata = 32'd21685;
			43852: outdata = 32'd21684;
			43853: outdata = 32'd21683;
			43854: outdata = 32'd21682;
			43855: outdata = 32'd21681;
			43856: outdata = 32'd21680;
			43857: outdata = 32'd21679;
			43858: outdata = 32'd21678;
			43859: outdata = 32'd21677;
			43860: outdata = 32'd21676;
			43861: outdata = 32'd21675;
			43862: outdata = 32'd21674;
			43863: outdata = 32'd21673;
			43864: outdata = 32'd21672;
			43865: outdata = 32'd21671;
			43866: outdata = 32'd21670;
			43867: outdata = 32'd21669;
			43868: outdata = 32'd21668;
			43869: outdata = 32'd21667;
			43870: outdata = 32'd21666;
			43871: outdata = 32'd21665;
			43872: outdata = 32'd21664;
			43873: outdata = 32'd21663;
			43874: outdata = 32'd21662;
			43875: outdata = 32'd21661;
			43876: outdata = 32'd21660;
			43877: outdata = 32'd21659;
			43878: outdata = 32'd21658;
			43879: outdata = 32'd21657;
			43880: outdata = 32'd21656;
			43881: outdata = 32'd21655;
			43882: outdata = 32'd21654;
			43883: outdata = 32'd21653;
			43884: outdata = 32'd21652;
			43885: outdata = 32'd21651;
			43886: outdata = 32'd21650;
			43887: outdata = 32'd21649;
			43888: outdata = 32'd21648;
			43889: outdata = 32'd21647;
			43890: outdata = 32'd21646;
			43891: outdata = 32'd21645;
			43892: outdata = 32'd21644;
			43893: outdata = 32'd21643;
			43894: outdata = 32'd21642;
			43895: outdata = 32'd21641;
			43896: outdata = 32'd21640;
			43897: outdata = 32'd21639;
			43898: outdata = 32'd21638;
			43899: outdata = 32'd21637;
			43900: outdata = 32'd21636;
			43901: outdata = 32'd21635;
			43902: outdata = 32'd21634;
			43903: outdata = 32'd21633;
			43904: outdata = 32'd21632;
			43905: outdata = 32'd21631;
			43906: outdata = 32'd21630;
			43907: outdata = 32'd21629;
			43908: outdata = 32'd21628;
			43909: outdata = 32'd21627;
			43910: outdata = 32'd21626;
			43911: outdata = 32'd21625;
			43912: outdata = 32'd21624;
			43913: outdata = 32'd21623;
			43914: outdata = 32'd21622;
			43915: outdata = 32'd21621;
			43916: outdata = 32'd21620;
			43917: outdata = 32'd21619;
			43918: outdata = 32'd21618;
			43919: outdata = 32'd21617;
			43920: outdata = 32'd21616;
			43921: outdata = 32'd21615;
			43922: outdata = 32'd21614;
			43923: outdata = 32'd21613;
			43924: outdata = 32'd21612;
			43925: outdata = 32'd21611;
			43926: outdata = 32'd21610;
			43927: outdata = 32'd21609;
			43928: outdata = 32'd21608;
			43929: outdata = 32'd21607;
			43930: outdata = 32'd21606;
			43931: outdata = 32'd21605;
			43932: outdata = 32'd21604;
			43933: outdata = 32'd21603;
			43934: outdata = 32'd21602;
			43935: outdata = 32'd21601;
			43936: outdata = 32'd21600;
			43937: outdata = 32'd21599;
			43938: outdata = 32'd21598;
			43939: outdata = 32'd21597;
			43940: outdata = 32'd21596;
			43941: outdata = 32'd21595;
			43942: outdata = 32'd21594;
			43943: outdata = 32'd21593;
			43944: outdata = 32'd21592;
			43945: outdata = 32'd21591;
			43946: outdata = 32'd21590;
			43947: outdata = 32'd21589;
			43948: outdata = 32'd21588;
			43949: outdata = 32'd21587;
			43950: outdata = 32'd21586;
			43951: outdata = 32'd21585;
			43952: outdata = 32'd21584;
			43953: outdata = 32'd21583;
			43954: outdata = 32'd21582;
			43955: outdata = 32'd21581;
			43956: outdata = 32'd21580;
			43957: outdata = 32'd21579;
			43958: outdata = 32'd21578;
			43959: outdata = 32'd21577;
			43960: outdata = 32'd21576;
			43961: outdata = 32'd21575;
			43962: outdata = 32'd21574;
			43963: outdata = 32'd21573;
			43964: outdata = 32'd21572;
			43965: outdata = 32'd21571;
			43966: outdata = 32'd21570;
			43967: outdata = 32'd21569;
			43968: outdata = 32'd21568;
			43969: outdata = 32'd21567;
			43970: outdata = 32'd21566;
			43971: outdata = 32'd21565;
			43972: outdata = 32'd21564;
			43973: outdata = 32'd21563;
			43974: outdata = 32'd21562;
			43975: outdata = 32'd21561;
			43976: outdata = 32'd21560;
			43977: outdata = 32'd21559;
			43978: outdata = 32'd21558;
			43979: outdata = 32'd21557;
			43980: outdata = 32'd21556;
			43981: outdata = 32'd21555;
			43982: outdata = 32'd21554;
			43983: outdata = 32'd21553;
			43984: outdata = 32'd21552;
			43985: outdata = 32'd21551;
			43986: outdata = 32'd21550;
			43987: outdata = 32'd21549;
			43988: outdata = 32'd21548;
			43989: outdata = 32'd21547;
			43990: outdata = 32'd21546;
			43991: outdata = 32'd21545;
			43992: outdata = 32'd21544;
			43993: outdata = 32'd21543;
			43994: outdata = 32'd21542;
			43995: outdata = 32'd21541;
			43996: outdata = 32'd21540;
			43997: outdata = 32'd21539;
			43998: outdata = 32'd21538;
			43999: outdata = 32'd21537;
			44000: outdata = 32'd21536;
			44001: outdata = 32'd21535;
			44002: outdata = 32'd21534;
			44003: outdata = 32'd21533;
			44004: outdata = 32'd21532;
			44005: outdata = 32'd21531;
			44006: outdata = 32'd21530;
			44007: outdata = 32'd21529;
			44008: outdata = 32'd21528;
			44009: outdata = 32'd21527;
			44010: outdata = 32'd21526;
			44011: outdata = 32'd21525;
			44012: outdata = 32'd21524;
			44013: outdata = 32'd21523;
			44014: outdata = 32'd21522;
			44015: outdata = 32'd21521;
			44016: outdata = 32'd21520;
			44017: outdata = 32'd21519;
			44018: outdata = 32'd21518;
			44019: outdata = 32'd21517;
			44020: outdata = 32'd21516;
			44021: outdata = 32'd21515;
			44022: outdata = 32'd21514;
			44023: outdata = 32'd21513;
			44024: outdata = 32'd21512;
			44025: outdata = 32'd21511;
			44026: outdata = 32'd21510;
			44027: outdata = 32'd21509;
			44028: outdata = 32'd21508;
			44029: outdata = 32'd21507;
			44030: outdata = 32'd21506;
			44031: outdata = 32'd21505;
			44032: outdata = 32'd21504;
			44033: outdata = 32'd21503;
			44034: outdata = 32'd21502;
			44035: outdata = 32'd21501;
			44036: outdata = 32'd21500;
			44037: outdata = 32'd21499;
			44038: outdata = 32'd21498;
			44039: outdata = 32'd21497;
			44040: outdata = 32'd21496;
			44041: outdata = 32'd21495;
			44042: outdata = 32'd21494;
			44043: outdata = 32'd21493;
			44044: outdata = 32'd21492;
			44045: outdata = 32'd21491;
			44046: outdata = 32'd21490;
			44047: outdata = 32'd21489;
			44048: outdata = 32'd21488;
			44049: outdata = 32'd21487;
			44050: outdata = 32'd21486;
			44051: outdata = 32'd21485;
			44052: outdata = 32'd21484;
			44053: outdata = 32'd21483;
			44054: outdata = 32'd21482;
			44055: outdata = 32'd21481;
			44056: outdata = 32'd21480;
			44057: outdata = 32'd21479;
			44058: outdata = 32'd21478;
			44059: outdata = 32'd21477;
			44060: outdata = 32'd21476;
			44061: outdata = 32'd21475;
			44062: outdata = 32'd21474;
			44063: outdata = 32'd21473;
			44064: outdata = 32'd21472;
			44065: outdata = 32'd21471;
			44066: outdata = 32'd21470;
			44067: outdata = 32'd21469;
			44068: outdata = 32'd21468;
			44069: outdata = 32'd21467;
			44070: outdata = 32'd21466;
			44071: outdata = 32'd21465;
			44072: outdata = 32'd21464;
			44073: outdata = 32'd21463;
			44074: outdata = 32'd21462;
			44075: outdata = 32'd21461;
			44076: outdata = 32'd21460;
			44077: outdata = 32'd21459;
			44078: outdata = 32'd21458;
			44079: outdata = 32'd21457;
			44080: outdata = 32'd21456;
			44081: outdata = 32'd21455;
			44082: outdata = 32'd21454;
			44083: outdata = 32'd21453;
			44084: outdata = 32'd21452;
			44085: outdata = 32'd21451;
			44086: outdata = 32'd21450;
			44087: outdata = 32'd21449;
			44088: outdata = 32'd21448;
			44089: outdata = 32'd21447;
			44090: outdata = 32'd21446;
			44091: outdata = 32'd21445;
			44092: outdata = 32'd21444;
			44093: outdata = 32'd21443;
			44094: outdata = 32'd21442;
			44095: outdata = 32'd21441;
			44096: outdata = 32'd21440;
			44097: outdata = 32'd21439;
			44098: outdata = 32'd21438;
			44099: outdata = 32'd21437;
			44100: outdata = 32'd21436;
			44101: outdata = 32'd21435;
			44102: outdata = 32'd21434;
			44103: outdata = 32'd21433;
			44104: outdata = 32'd21432;
			44105: outdata = 32'd21431;
			44106: outdata = 32'd21430;
			44107: outdata = 32'd21429;
			44108: outdata = 32'd21428;
			44109: outdata = 32'd21427;
			44110: outdata = 32'd21426;
			44111: outdata = 32'd21425;
			44112: outdata = 32'd21424;
			44113: outdata = 32'd21423;
			44114: outdata = 32'd21422;
			44115: outdata = 32'd21421;
			44116: outdata = 32'd21420;
			44117: outdata = 32'd21419;
			44118: outdata = 32'd21418;
			44119: outdata = 32'd21417;
			44120: outdata = 32'd21416;
			44121: outdata = 32'd21415;
			44122: outdata = 32'd21414;
			44123: outdata = 32'd21413;
			44124: outdata = 32'd21412;
			44125: outdata = 32'd21411;
			44126: outdata = 32'd21410;
			44127: outdata = 32'd21409;
			44128: outdata = 32'd21408;
			44129: outdata = 32'd21407;
			44130: outdata = 32'd21406;
			44131: outdata = 32'd21405;
			44132: outdata = 32'd21404;
			44133: outdata = 32'd21403;
			44134: outdata = 32'd21402;
			44135: outdata = 32'd21401;
			44136: outdata = 32'd21400;
			44137: outdata = 32'd21399;
			44138: outdata = 32'd21398;
			44139: outdata = 32'd21397;
			44140: outdata = 32'd21396;
			44141: outdata = 32'd21395;
			44142: outdata = 32'd21394;
			44143: outdata = 32'd21393;
			44144: outdata = 32'd21392;
			44145: outdata = 32'd21391;
			44146: outdata = 32'd21390;
			44147: outdata = 32'd21389;
			44148: outdata = 32'd21388;
			44149: outdata = 32'd21387;
			44150: outdata = 32'd21386;
			44151: outdata = 32'd21385;
			44152: outdata = 32'd21384;
			44153: outdata = 32'd21383;
			44154: outdata = 32'd21382;
			44155: outdata = 32'd21381;
			44156: outdata = 32'd21380;
			44157: outdata = 32'd21379;
			44158: outdata = 32'd21378;
			44159: outdata = 32'd21377;
			44160: outdata = 32'd21376;
			44161: outdata = 32'd21375;
			44162: outdata = 32'd21374;
			44163: outdata = 32'd21373;
			44164: outdata = 32'd21372;
			44165: outdata = 32'd21371;
			44166: outdata = 32'd21370;
			44167: outdata = 32'd21369;
			44168: outdata = 32'd21368;
			44169: outdata = 32'd21367;
			44170: outdata = 32'd21366;
			44171: outdata = 32'd21365;
			44172: outdata = 32'd21364;
			44173: outdata = 32'd21363;
			44174: outdata = 32'd21362;
			44175: outdata = 32'd21361;
			44176: outdata = 32'd21360;
			44177: outdata = 32'd21359;
			44178: outdata = 32'd21358;
			44179: outdata = 32'd21357;
			44180: outdata = 32'd21356;
			44181: outdata = 32'd21355;
			44182: outdata = 32'd21354;
			44183: outdata = 32'd21353;
			44184: outdata = 32'd21352;
			44185: outdata = 32'd21351;
			44186: outdata = 32'd21350;
			44187: outdata = 32'd21349;
			44188: outdata = 32'd21348;
			44189: outdata = 32'd21347;
			44190: outdata = 32'd21346;
			44191: outdata = 32'd21345;
			44192: outdata = 32'd21344;
			44193: outdata = 32'd21343;
			44194: outdata = 32'd21342;
			44195: outdata = 32'd21341;
			44196: outdata = 32'd21340;
			44197: outdata = 32'd21339;
			44198: outdata = 32'd21338;
			44199: outdata = 32'd21337;
			44200: outdata = 32'd21336;
			44201: outdata = 32'd21335;
			44202: outdata = 32'd21334;
			44203: outdata = 32'd21333;
			44204: outdata = 32'd21332;
			44205: outdata = 32'd21331;
			44206: outdata = 32'd21330;
			44207: outdata = 32'd21329;
			44208: outdata = 32'd21328;
			44209: outdata = 32'd21327;
			44210: outdata = 32'd21326;
			44211: outdata = 32'd21325;
			44212: outdata = 32'd21324;
			44213: outdata = 32'd21323;
			44214: outdata = 32'd21322;
			44215: outdata = 32'd21321;
			44216: outdata = 32'd21320;
			44217: outdata = 32'd21319;
			44218: outdata = 32'd21318;
			44219: outdata = 32'd21317;
			44220: outdata = 32'd21316;
			44221: outdata = 32'd21315;
			44222: outdata = 32'd21314;
			44223: outdata = 32'd21313;
			44224: outdata = 32'd21312;
			44225: outdata = 32'd21311;
			44226: outdata = 32'd21310;
			44227: outdata = 32'd21309;
			44228: outdata = 32'd21308;
			44229: outdata = 32'd21307;
			44230: outdata = 32'd21306;
			44231: outdata = 32'd21305;
			44232: outdata = 32'd21304;
			44233: outdata = 32'd21303;
			44234: outdata = 32'd21302;
			44235: outdata = 32'd21301;
			44236: outdata = 32'd21300;
			44237: outdata = 32'd21299;
			44238: outdata = 32'd21298;
			44239: outdata = 32'd21297;
			44240: outdata = 32'd21296;
			44241: outdata = 32'd21295;
			44242: outdata = 32'd21294;
			44243: outdata = 32'd21293;
			44244: outdata = 32'd21292;
			44245: outdata = 32'd21291;
			44246: outdata = 32'd21290;
			44247: outdata = 32'd21289;
			44248: outdata = 32'd21288;
			44249: outdata = 32'd21287;
			44250: outdata = 32'd21286;
			44251: outdata = 32'd21285;
			44252: outdata = 32'd21284;
			44253: outdata = 32'd21283;
			44254: outdata = 32'd21282;
			44255: outdata = 32'd21281;
			44256: outdata = 32'd21280;
			44257: outdata = 32'd21279;
			44258: outdata = 32'd21278;
			44259: outdata = 32'd21277;
			44260: outdata = 32'd21276;
			44261: outdata = 32'd21275;
			44262: outdata = 32'd21274;
			44263: outdata = 32'd21273;
			44264: outdata = 32'd21272;
			44265: outdata = 32'd21271;
			44266: outdata = 32'd21270;
			44267: outdata = 32'd21269;
			44268: outdata = 32'd21268;
			44269: outdata = 32'd21267;
			44270: outdata = 32'd21266;
			44271: outdata = 32'd21265;
			44272: outdata = 32'd21264;
			44273: outdata = 32'd21263;
			44274: outdata = 32'd21262;
			44275: outdata = 32'd21261;
			44276: outdata = 32'd21260;
			44277: outdata = 32'd21259;
			44278: outdata = 32'd21258;
			44279: outdata = 32'd21257;
			44280: outdata = 32'd21256;
			44281: outdata = 32'd21255;
			44282: outdata = 32'd21254;
			44283: outdata = 32'd21253;
			44284: outdata = 32'd21252;
			44285: outdata = 32'd21251;
			44286: outdata = 32'd21250;
			44287: outdata = 32'd21249;
			44288: outdata = 32'd21248;
			44289: outdata = 32'd21247;
			44290: outdata = 32'd21246;
			44291: outdata = 32'd21245;
			44292: outdata = 32'd21244;
			44293: outdata = 32'd21243;
			44294: outdata = 32'd21242;
			44295: outdata = 32'd21241;
			44296: outdata = 32'd21240;
			44297: outdata = 32'd21239;
			44298: outdata = 32'd21238;
			44299: outdata = 32'd21237;
			44300: outdata = 32'd21236;
			44301: outdata = 32'd21235;
			44302: outdata = 32'd21234;
			44303: outdata = 32'd21233;
			44304: outdata = 32'd21232;
			44305: outdata = 32'd21231;
			44306: outdata = 32'd21230;
			44307: outdata = 32'd21229;
			44308: outdata = 32'd21228;
			44309: outdata = 32'd21227;
			44310: outdata = 32'd21226;
			44311: outdata = 32'd21225;
			44312: outdata = 32'd21224;
			44313: outdata = 32'd21223;
			44314: outdata = 32'd21222;
			44315: outdata = 32'd21221;
			44316: outdata = 32'd21220;
			44317: outdata = 32'd21219;
			44318: outdata = 32'd21218;
			44319: outdata = 32'd21217;
			44320: outdata = 32'd21216;
			44321: outdata = 32'd21215;
			44322: outdata = 32'd21214;
			44323: outdata = 32'd21213;
			44324: outdata = 32'd21212;
			44325: outdata = 32'd21211;
			44326: outdata = 32'd21210;
			44327: outdata = 32'd21209;
			44328: outdata = 32'd21208;
			44329: outdata = 32'd21207;
			44330: outdata = 32'd21206;
			44331: outdata = 32'd21205;
			44332: outdata = 32'd21204;
			44333: outdata = 32'd21203;
			44334: outdata = 32'd21202;
			44335: outdata = 32'd21201;
			44336: outdata = 32'd21200;
			44337: outdata = 32'd21199;
			44338: outdata = 32'd21198;
			44339: outdata = 32'd21197;
			44340: outdata = 32'd21196;
			44341: outdata = 32'd21195;
			44342: outdata = 32'd21194;
			44343: outdata = 32'd21193;
			44344: outdata = 32'd21192;
			44345: outdata = 32'd21191;
			44346: outdata = 32'd21190;
			44347: outdata = 32'd21189;
			44348: outdata = 32'd21188;
			44349: outdata = 32'd21187;
			44350: outdata = 32'd21186;
			44351: outdata = 32'd21185;
			44352: outdata = 32'd21184;
			44353: outdata = 32'd21183;
			44354: outdata = 32'd21182;
			44355: outdata = 32'd21181;
			44356: outdata = 32'd21180;
			44357: outdata = 32'd21179;
			44358: outdata = 32'd21178;
			44359: outdata = 32'd21177;
			44360: outdata = 32'd21176;
			44361: outdata = 32'd21175;
			44362: outdata = 32'd21174;
			44363: outdata = 32'd21173;
			44364: outdata = 32'd21172;
			44365: outdata = 32'd21171;
			44366: outdata = 32'd21170;
			44367: outdata = 32'd21169;
			44368: outdata = 32'd21168;
			44369: outdata = 32'd21167;
			44370: outdata = 32'd21166;
			44371: outdata = 32'd21165;
			44372: outdata = 32'd21164;
			44373: outdata = 32'd21163;
			44374: outdata = 32'd21162;
			44375: outdata = 32'd21161;
			44376: outdata = 32'd21160;
			44377: outdata = 32'd21159;
			44378: outdata = 32'd21158;
			44379: outdata = 32'd21157;
			44380: outdata = 32'd21156;
			44381: outdata = 32'd21155;
			44382: outdata = 32'd21154;
			44383: outdata = 32'd21153;
			44384: outdata = 32'd21152;
			44385: outdata = 32'd21151;
			44386: outdata = 32'd21150;
			44387: outdata = 32'd21149;
			44388: outdata = 32'd21148;
			44389: outdata = 32'd21147;
			44390: outdata = 32'd21146;
			44391: outdata = 32'd21145;
			44392: outdata = 32'd21144;
			44393: outdata = 32'd21143;
			44394: outdata = 32'd21142;
			44395: outdata = 32'd21141;
			44396: outdata = 32'd21140;
			44397: outdata = 32'd21139;
			44398: outdata = 32'd21138;
			44399: outdata = 32'd21137;
			44400: outdata = 32'd21136;
			44401: outdata = 32'd21135;
			44402: outdata = 32'd21134;
			44403: outdata = 32'd21133;
			44404: outdata = 32'd21132;
			44405: outdata = 32'd21131;
			44406: outdata = 32'd21130;
			44407: outdata = 32'd21129;
			44408: outdata = 32'd21128;
			44409: outdata = 32'd21127;
			44410: outdata = 32'd21126;
			44411: outdata = 32'd21125;
			44412: outdata = 32'd21124;
			44413: outdata = 32'd21123;
			44414: outdata = 32'd21122;
			44415: outdata = 32'd21121;
			44416: outdata = 32'd21120;
			44417: outdata = 32'd21119;
			44418: outdata = 32'd21118;
			44419: outdata = 32'd21117;
			44420: outdata = 32'd21116;
			44421: outdata = 32'd21115;
			44422: outdata = 32'd21114;
			44423: outdata = 32'd21113;
			44424: outdata = 32'd21112;
			44425: outdata = 32'd21111;
			44426: outdata = 32'd21110;
			44427: outdata = 32'd21109;
			44428: outdata = 32'd21108;
			44429: outdata = 32'd21107;
			44430: outdata = 32'd21106;
			44431: outdata = 32'd21105;
			44432: outdata = 32'd21104;
			44433: outdata = 32'd21103;
			44434: outdata = 32'd21102;
			44435: outdata = 32'd21101;
			44436: outdata = 32'd21100;
			44437: outdata = 32'd21099;
			44438: outdata = 32'd21098;
			44439: outdata = 32'd21097;
			44440: outdata = 32'd21096;
			44441: outdata = 32'd21095;
			44442: outdata = 32'd21094;
			44443: outdata = 32'd21093;
			44444: outdata = 32'd21092;
			44445: outdata = 32'd21091;
			44446: outdata = 32'd21090;
			44447: outdata = 32'd21089;
			44448: outdata = 32'd21088;
			44449: outdata = 32'd21087;
			44450: outdata = 32'd21086;
			44451: outdata = 32'd21085;
			44452: outdata = 32'd21084;
			44453: outdata = 32'd21083;
			44454: outdata = 32'd21082;
			44455: outdata = 32'd21081;
			44456: outdata = 32'd21080;
			44457: outdata = 32'd21079;
			44458: outdata = 32'd21078;
			44459: outdata = 32'd21077;
			44460: outdata = 32'd21076;
			44461: outdata = 32'd21075;
			44462: outdata = 32'd21074;
			44463: outdata = 32'd21073;
			44464: outdata = 32'd21072;
			44465: outdata = 32'd21071;
			44466: outdata = 32'd21070;
			44467: outdata = 32'd21069;
			44468: outdata = 32'd21068;
			44469: outdata = 32'd21067;
			44470: outdata = 32'd21066;
			44471: outdata = 32'd21065;
			44472: outdata = 32'd21064;
			44473: outdata = 32'd21063;
			44474: outdata = 32'd21062;
			44475: outdata = 32'd21061;
			44476: outdata = 32'd21060;
			44477: outdata = 32'd21059;
			44478: outdata = 32'd21058;
			44479: outdata = 32'd21057;
			44480: outdata = 32'd21056;
			44481: outdata = 32'd21055;
			44482: outdata = 32'd21054;
			44483: outdata = 32'd21053;
			44484: outdata = 32'd21052;
			44485: outdata = 32'd21051;
			44486: outdata = 32'd21050;
			44487: outdata = 32'd21049;
			44488: outdata = 32'd21048;
			44489: outdata = 32'd21047;
			44490: outdata = 32'd21046;
			44491: outdata = 32'd21045;
			44492: outdata = 32'd21044;
			44493: outdata = 32'd21043;
			44494: outdata = 32'd21042;
			44495: outdata = 32'd21041;
			44496: outdata = 32'd21040;
			44497: outdata = 32'd21039;
			44498: outdata = 32'd21038;
			44499: outdata = 32'd21037;
			44500: outdata = 32'd21036;
			44501: outdata = 32'd21035;
			44502: outdata = 32'd21034;
			44503: outdata = 32'd21033;
			44504: outdata = 32'd21032;
			44505: outdata = 32'd21031;
			44506: outdata = 32'd21030;
			44507: outdata = 32'd21029;
			44508: outdata = 32'd21028;
			44509: outdata = 32'd21027;
			44510: outdata = 32'd21026;
			44511: outdata = 32'd21025;
			44512: outdata = 32'd21024;
			44513: outdata = 32'd21023;
			44514: outdata = 32'd21022;
			44515: outdata = 32'd21021;
			44516: outdata = 32'd21020;
			44517: outdata = 32'd21019;
			44518: outdata = 32'd21018;
			44519: outdata = 32'd21017;
			44520: outdata = 32'd21016;
			44521: outdata = 32'd21015;
			44522: outdata = 32'd21014;
			44523: outdata = 32'd21013;
			44524: outdata = 32'd21012;
			44525: outdata = 32'd21011;
			44526: outdata = 32'd21010;
			44527: outdata = 32'd21009;
			44528: outdata = 32'd21008;
			44529: outdata = 32'd21007;
			44530: outdata = 32'd21006;
			44531: outdata = 32'd21005;
			44532: outdata = 32'd21004;
			44533: outdata = 32'd21003;
			44534: outdata = 32'd21002;
			44535: outdata = 32'd21001;
			44536: outdata = 32'd21000;
			44537: outdata = 32'd20999;
			44538: outdata = 32'd20998;
			44539: outdata = 32'd20997;
			44540: outdata = 32'd20996;
			44541: outdata = 32'd20995;
			44542: outdata = 32'd20994;
			44543: outdata = 32'd20993;
			44544: outdata = 32'd20992;
			44545: outdata = 32'd20991;
			44546: outdata = 32'd20990;
			44547: outdata = 32'd20989;
			44548: outdata = 32'd20988;
			44549: outdata = 32'd20987;
			44550: outdata = 32'd20986;
			44551: outdata = 32'd20985;
			44552: outdata = 32'd20984;
			44553: outdata = 32'd20983;
			44554: outdata = 32'd20982;
			44555: outdata = 32'd20981;
			44556: outdata = 32'd20980;
			44557: outdata = 32'd20979;
			44558: outdata = 32'd20978;
			44559: outdata = 32'd20977;
			44560: outdata = 32'd20976;
			44561: outdata = 32'd20975;
			44562: outdata = 32'd20974;
			44563: outdata = 32'd20973;
			44564: outdata = 32'd20972;
			44565: outdata = 32'd20971;
			44566: outdata = 32'd20970;
			44567: outdata = 32'd20969;
			44568: outdata = 32'd20968;
			44569: outdata = 32'd20967;
			44570: outdata = 32'd20966;
			44571: outdata = 32'd20965;
			44572: outdata = 32'd20964;
			44573: outdata = 32'd20963;
			44574: outdata = 32'd20962;
			44575: outdata = 32'd20961;
			44576: outdata = 32'd20960;
			44577: outdata = 32'd20959;
			44578: outdata = 32'd20958;
			44579: outdata = 32'd20957;
			44580: outdata = 32'd20956;
			44581: outdata = 32'd20955;
			44582: outdata = 32'd20954;
			44583: outdata = 32'd20953;
			44584: outdata = 32'd20952;
			44585: outdata = 32'd20951;
			44586: outdata = 32'd20950;
			44587: outdata = 32'd20949;
			44588: outdata = 32'd20948;
			44589: outdata = 32'd20947;
			44590: outdata = 32'd20946;
			44591: outdata = 32'd20945;
			44592: outdata = 32'd20944;
			44593: outdata = 32'd20943;
			44594: outdata = 32'd20942;
			44595: outdata = 32'd20941;
			44596: outdata = 32'd20940;
			44597: outdata = 32'd20939;
			44598: outdata = 32'd20938;
			44599: outdata = 32'd20937;
			44600: outdata = 32'd20936;
			44601: outdata = 32'd20935;
			44602: outdata = 32'd20934;
			44603: outdata = 32'd20933;
			44604: outdata = 32'd20932;
			44605: outdata = 32'd20931;
			44606: outdata = 32'd20930;
			44607: outdata = 32'd20929;
			44608: outdata = 32'd20928;
			44609: outdata = 32'd20927;
			44610: outdata = 32'd20926;
			44611: outdata = 32'd20925;
			44612: outdata = 32'd20924;
			44613: outdata = 32'd20923;
			44614: outdata = 32'd20922;
			44615: outdata = 32'd20921;
			44616: outdata = 32'd20920;
			44617: outdata = 32'd20919;
			44618: outdata = 32'd20918;
			44619: outdata = 32'd20917;
			44620: outdata = 32'd20916;
			44621: outdata = 32'd20915;
			44622: outdata = 32'd20914;
			44623: outdata = 32'd20913;
			44624: outdata = 32'd20912;
			44625: outdata = 32'd20911;
			44626: outdata = 32'd20910;
			44627: outdata = 32'd20909;
			44628: outdata = 32'd20908;
			44629: outdata = 32'd20907;
			44630: outdata = 32'd20906;
			44631: outdata = 32'd20905;
			44632: outdata = 32'd20904;
			44633: outdata = 32'd20903;
			44634: outdata = 32'd20902;
			44635: outdata = 32'd20901;
			44636: outdata = 32'd20900;
			44637: outdata = 32'd20899;
			44638: outdata = 32'd20898;
			44639: outdata = 32'd20897;
			44640: outdata = 32'd20896;
			44641: outdata = 32'd20895;
			44642: outdata = 32'd20894;
			44643: outdata = 32'd20893;
			44644: outdata = 32'd20892;
			44645: outdata = 32'd20891;
			44646: outdata = 32'd20890;
			44647: outdata = 32'd20889;
			44648: outdata = 32'd20888;
			44649: outdata = 32'd20887;
			44650: outdata = 32'd20886;
			44651: outdata = 32'd20885;
			44652: outdata = 32'd20884;
			44653: outdata = 32'd20883;
			44654: outdata = 32'd20882;
			44655: outdata = 32'd20881;
			44656: outdata = 32'd20880;
			44657: outdata = 32'd20879;
			44658: outdata = 32'd20878;
			44659: outdata = 32'd20877;
			44660: outdata = 32'd20876;
			44661: outdata = 32'd20875;
			44662: outdata = 32'd20874;
			44663: outdata = 32'd20873;
			44664: outdata = 32'd20872;
			44665: outdata = 32'd20871;
			44666: outdata = 32'd20870;
			44667: outdata = 32'd20869;
			44668: outdata = 32'd20868;
			44669: outdata = 32'd20867;
			44670: outdata = 32'd20866;
			44671: outdata = 32'd20865;
			44672: outdata = 32'd20864;
			44673: outdata = 32'd20863;
			44674: outdata = 32'd20862;
			44675: outdata = 32'd20861;
			44676: outdata = 32'd20860;
			44677: outdata = 32'd20859;
			44678: outdata = 32'd20858;
			44679: outdata = 32'd20857;
			44680: outdata = 32'd20856;
			44681: outdata = 32'd20855;
			44682: outdata = 32'd20854;
			44683: outdata = 32'd20853;
			44684: outdata = 32'd20852;
			44685: outdata = 32'd20851;
			44686: outdata = 32'd20850;
			44687: outdata = 32'd20849;
			44688: outdata = 32'd20848;
			44689: outdata = 32'd20847;
			44690: outdata = 32'd20846;
			44691: outdata = 32'd20845;
			44692: outdata = 32'd20844;
			44693: outdata = 32'd20843;
			44694: outdata = 32'd20842;
			44695: outdata = 32'd20841;
			44696: outdata = 32'd20840;
			44697: outdata = 32'd20839;
			44698: outdata = 32'd20838;
			44699: outdata = 32'd20837;
			44700: outdata = 32'd20836;
			44701: outdata = 32'd20835;
			44702: outdata = 32'd20834;
			44703: outdata = 32'd20833;
			44704: outdata = 32'd20832;
			44705: outdata = 32'd20831;
			44706: outdata = 32'd20830;
			44707: outdata = 32'd20829;
			44708: outdata = 32'd20828;
			44709: outdata = 32'd20827;
			44710: outdata = 32'd20826;
			44711: outdata = 32'd20825;
			44712: outdata = 32'd20824;
			44713: outdata = 32'd20823;
			44714: outdata = 32'd20822;
			44715: outdata = 32'd20821;
			44716: outdata = 32'd20820;
			44717: outdata = 32'd20819;
			44718: outdata = 32'd20818;
			44719: outdata = 32'd20817;
			44720: outdata = 32'd20816;
			44721: outdata = 32'd20815;
			44722: outdata = 32'd20814;
			44723: outdata = 32'd20813;
			44724: outdata = 32'd20812;
			44725: outdata = 32'd20811;
			44726: outdata = 32'd20810;
			44727: outdata = 32'd20809;
			44728: outdata = 32'd20808;
			44729: outdata = 32'd20807;
			44730: outdata = 32'd20806;
			44731: outdata = 32'd20805;
			44732: outdata = 32'd20804;
			44733: outdata = 32'd20803;
			44734: outdata = 32'd20802;
			44735: outdata = 32'd20801;
			44736: outdata = 32'd20800;
			44737: outdata = 32'd20799;
			44738: outdata = 32'd20798;
			44739: outdata = 32'd20797;
			44740: outdata = 32'd20796;
			44741: outdata = 32'd20795;
			44742: outdata = 32'd20794;
			44743: outdata = 32'd20793;
			44744: outdata = 32'd20792;
			44745: outdata = 32'd20791;
			44746: outdata = 32'd20790;
			44747: outdata = 32'd20789;
			44748: outdata = 32'd20788;
			44749: outdata = 32'd20787;
			44750: outdata = 32'd20786;
			44751: outdata = 32'd20785;
			44752: outdata = 32'd20784;
			44753: outdata = 32'd20783;
			44754: outdata = 32'd20782;
			44755: outdata = 32'd20781;
			44756: outdata = 32'd20780;
			44757: outdata = 32'd20779;
			44758: outdata = 32'd20778;
			44759: outdata = 32'd20777;
			44760: outdata = 32'd20776;
			44761: outdata = 32'd20775;
			44762: outdata = 32'd20774;
			44763: outdata = 32'd20773;
			44764: outdata = 32'd20772;
			44765: outdata = 32'd20771;
			44766: outdata = 32'd20770;
			44767: outdata = 32'd20769;
			44768: outdata = 32'd20768;
			44769: outdata = 32'd20767;
			44770: outdata = 32'd20766;
			44771: outdata = 32'd20765;
			44772: outdata = 32'd20764;
			44773: outdata = 32'd20763;
			44774: outdata = 32'd20762;
			44775: outdata = 32'd20761;
			44776: outdata = 32'd20760;
			44777: outdata = 32'd20759;
			44778: outdata = 32'd20758;
			44779: outdata = 32'd20757;
			44780: outdata = 32'd20756;
			44781: outdata = 32'd20755;
			44782: outdata = 32'd20754;
			44783: outdata = 32'd20753;
			44784: outdata = 32'd20752;
			44785: outdata = 32'd20751;
			44786: outdata = 32'd20750;
			44787: outdata = 32'd20749;
			44788: outdata = 32'd20748;
			44789: outdata = 32'd20747;
			44790: outdata = 32'd20746;
			44791: outdata = 32'd20745;
			44792: outdata = 32'd20744;
			44793: outdata = 32'd20743;
			44794: outdata = 32'd20742;
			44795: outdata = 32'd20741;
			44796: outdata = 32'd20740;
			44797: outdata = 32'd20739;
			44798: outdata = 32'd20738;
			44799: outdata = 32'd20737;
			44800: outdata = 32'd20736;
			44801: outdata = 32'd20735;
			44802: outdata = 32'd20734;
			44803: outdata = 32'd20733;
			44804: outdata = 32'd20732;
			44805: outdata = 32'd20731;
			44806: outdata = 32'd20730;
			44807: outdata = 32'd20729;
			44808: outdata = 32'd20728;
			44809: outdata = 32'd20727;
			44810: outdata = 32'd20726;
			44811: outdata = 32'd20725;
			44812: outdata = 32'd20724;
			44813: outdata = 32'd20723;
			44814: outdata = 32'd20722;
			44815: outdata = 32'd20721;
			44816: outdata = 32'd20720;
			44817: outdata = 32'd20719;
			44818: outdata = 32'd20718;
			44819: outdata = 32'd20717;
			44820: outdata = 32'd20716;
			44821: outdata = 32'd20715;
			44822: outdata = 32'd20714;
			44823: outdata = 32'd20713;
			44824: outdata = 32'd20712;
			44825: outdata = 32'd20711;
			44826: outdata = 32'd20710;
			44827: outdata = 32'd20709;
			44828: outdata = 32'd20708;
			44829: outdata = 32'd20707;
			44830: outdata = 32'd20706;
			44831: outdata = 32'd20705;
			44832: outdata = 32'd20704;
			44833: outdata = 32'd20703;
			44834: outdata = 32'd20702;
			44835: outdata = 32'd20701;
			44836: outdata = 32'd20700;
			44837: outdata = 32'd20699;
			44838: outdata = 32'd20698;
			44839: outdata = 32'd20697;
			44840: outdata = 32'd20696;
			44841: outdata = 32'd20695;
			44842: outdata = 32'd20694;
			44843: outdata = 32'd20693;
			44844: outdata = 32'd20692;
			44845: outdata = 32'd20691;
			44846: outdata = 32'd20690;
			44847: outdata = 32'd20689;
			44848: outdata = 32'd20688;
			44849: outdata = 32'd20687;
			44850: outdata = 32'd20686;
			44851: outdata = 32'd20685;
			44852: outdata = 32'd20684;
			44853: outdata = 32'd20683;
			44854: outdata = 32'd20682;
			44855: outdata = 32'd20681;
			44856: outdata = 32'd20680;
			44857: outdata = 32'd20679;
			44858: outdata = 32'd20678;
			44859: outdata = 32'd20677;
			44860: outdata = 32'd20676;
			44861: outdata = 32'd20675;
			44862: outdata = 32'd20674;
			44863: outdata = 32'd20673;
			44864: outdata = 32'd20672;
			44865: outdata = 32'd20671;
			44866: outdata = 32'd20670;
			44867: outdata = 32'd20669;
			44868: outdata = 32'd20668;
			44869: outdata = 32'd20667;
			44870: outdata = 32'd20666;
			44871: outdata = 32'd20665;
			44872: outdata = 32'd20664;
			44873: outdata = 32'd20663;
			44874: outdata = 32'd20662;
			44875: outdata = 32'd20661;
			44876: outdata = 32'd20660;
			44877: outdata = 32'd20659;
			44878: outdata = 32'd20658;
			44879: outdata = 32'd20657;
			44880: outdata = 32'd20656;
			44881: outdata = 32'd20655;
			44882: outdata = 32'd20654;
			44883: outdata = 32'd20653;
			44884: outdata = 32'd20652;
			44885: outdata = 32'd20651;
			44886: outdata = 32'd20650;
			44887: outdata = 32'd20649;
			44888: outdata = 32'd20648;
			44889: outdata = 32'd20647;
			44890: outdata = 32'd20646;
			44891: outdata = 32'd20645;
			44892: outdata = 32'd20644;
			44893: outdata = 32'd20643;
			44894: outdata = 32'd20642;
			44895: outdata = 32'd20641;
			44896: outdata = 32'd20640;
			44897: outdata = 32'd20639;
			44898: outdata = 32'd20638;
			44899: outdata = 32'd20637;
			44900: outdata = 32'd20636;
			44901: outdata = 32'd20635;
			44902: outdata = 32'd20634;
			44903: outdata = 32'd20633;
			44904: outdata = 32'd20632;
			44905: outdata = 32'd20631;
			44906: outdata = 32'd20630;
			44907: outdata = 32'd20629;
			44908: outdata = 32'd20628;
			44909: outdata = 32'd20627;
			44910: outdata = 32'd20626;
			44911: outdata = 32'd20625;
			44912: outdata = 32'd20624;
			44913: outdata = 32'd20623;
			44914: outdata = 32'd20622;
			44915: outdata = 32'd20621;
			44916: outdata = 32'd20620;
			44917: outdata = 32'd20619;
			44918: outdata = 32'd20618;
			44919: outdata = 32'd20617;
			44920: outdata = 32'd20616;
			44921: outdata = 32'd20615;
			44922: outdata = 32'd20614;
			44923: outdata = 32'd20613;
			44924: outdata = 32'd20612;
			44925: outdata = 32'd20611;
			44926: outdata = 32'd20610;
			44927: outdata = 32'd20609;
			44928: outdata = 32'd20608;
			44929: outdata = 32'd20607;
			44930: outdata = 32'd20606;
			44931: outdata = 32'd20605;
			44932: outdata = 32'd20604;
			44933: outdata = 32'd20603;
			44934: outdata = 32'd20602;
			44935: outdata = 32'd20601;
			44936: outdata = 32'd20600;
			44937: outdata = 32'd20599;
			44938: outdata = 32'd20598;
			44939: outdata = 32'd20597;
			44940: outdata = 32'd20596;
			44941: outdata = 32'd20595;
			44942: outdata = 32'd20594;
			44943: outdata = 32'd20593;
			44944: outdata = 32'd20592;
			44945: outdata = 32'd20591;
			44946: outdata = 32'd20590;
			44947: outdata = 32'd20589;
			44948: outdata = 32'd20588;
			44949: outdata = 32'd20587;
			44950: outdata = 32'd20586;
			44951: outdata = 32'd20585;
			44952: outdata = 32'd20584;
			44953: outdata = 32'd20583;
			44954: outdata = 32'd20582;
			44955: outdata = 32'd20581;
			44956: outdata = 32'd20580;
			44957: outdata = 32'd20579;
			44958: outdata = 32'd20578;
			44959: outdata = 32'd20577;
			44960: outdata = 32'd20576;
			44961: outdata = 32'd20575;
			44962: outdata = 32'd20574;
			44963: outdata = 32'd20573;
			44964: outdata = 32'd20572;
			44965: outdata = 32'd20571;
			44966: outdata = 32'd20570;
			44967: outdata = 32'd20569;
			44968: outdata = 32'd20568;
			44969: outdata = 32'd20567;
			44970: outdata = 32'd20566;
			44971: outdata = 32'd20565;
			44972: outdata = 32'd20564;
			44973: outdata = 32'd20563;
			44974: outdata = 32'd20562;
			44975: outdata = 32'd20561;
			44976: outdata = 32'd20560;
			44977: outdata = 32'd20559;
			44978: outdata = 32'd20558;
			44979: outdata = 32'd20557;
			44980: outdata = 32'd20556;
			44981: outdata = 32'd20555;
			44982: outdata = 32'd20554;
			44983: outdata = 32'd20553;
			44984: outdata = 32'd20552;
			44985: outdata = 32'd20551;
			44986: outdata = 32'd20550;
			44987: outdata = 32'd20549;
			44988: outdata = 32'd20548;
			44989: outdata = 32'd20547;
			44990: outdata = 32'd20546;
			44991: outdata = 32'd20545;
			44992: outdata = 32'd20544;
			44993: outdata = 32'd20543;
			44994: outdata = 32'd20542;
			44995: outdata = 32'd20541;
			44996: outdata = 32'd20540;
			44997: outdata = 32'd20539;
			44998: outdata = 32'd20538;
			44999: outdata = 32'd20537;
			45000: outdata = 32'd20536;
			45001: outdata = 32'd20535;
			45002: outdata = 32'd20534;
			45003: outdata = 32'd20533;
			45004: outdata = 32'd20532;
			45005: outdata = 32'd20531;
			45006: outdata = 32'd20530;
			45007: outdata = 32'd20529;
			45008: outdata = 32'd20528;
			45009: outdata = 32'd20527;
			45010: outdata = 32'd20526;
			45011: outdata = 32'd20525;
			45012: outdata = 32'd20524;
			45013: outdata = 32'd20523;
			45014: outdata = 32'd20522;
			45015: outdata = 32'd20521;
			45016: outdata = 32'd20520;
			45017: outdata = 32'd20519;
			45018: outdata = 32'd20518;
			45019: outdata = 32'd20517;
			45020: outdata = 32'd20516;
			45021: outdata = 32'd20515;
			45022: outdata = 32'd20514;
			45023: outdata = 32'd20513;
			45024: outdata = 32'd20512;
			45025: outdata = 32'd20511;
			45026: outdata = 32'd20510;
			45027: outdata = 32'd20509;
			45028: outdata = 32'd20508;
			45029: outdata = 32'd20507;
			45030: outdata = 32'd20506;
			45031: outdata = 32'd20505;
			45032: outdata = 32'd20504;
			45033: outdata = 32'd20503;
			45034: outdata = 32'd20502;
			45035: outdata = 32'd20501;
			45036: outdata = 32'd20500;
			45037: outdata = 32'd20499;
			45038: outdata = 32'd20498;
			45039: outdata = 32'd20497;
			45040: outdata = 32'd20496;
			45041: outdata = 32'd20495;
			45042: outdata = 32'd20494;
			45043: outdata = 32'd20493;
			45044: outdata = 32'd20492;
			45045: outdata = 32'd20491;
			45046: outdata = 32'd20490;
			45047: outdata = 32'd20489;
			45048: outdata = 32'd20488;
			45049: outdata = 32'd20487;
			45050: outdata = 32'd20486;
			45051: outdata = 32'd20485;
			45052: outdata = 32'd20484;
			45053: outdata = 32'd20483;
			45054: outdata = 32'd20482;
			45055: outdata = 32'd20481;
			45056: outdata = 32'd20480;
			45057: outdata = 32'd20479;
			45058: outdata = 32'd20478;
			45059: outdata = 32'd20477;
			45060: outdata = 32'd20476;
			45061: outdata = 32'd20475;
			45062: outdata = 32'd20474;
			45063: outdata = 32'd20473;
			45064: outdata = 32'd20472;
			45065: outdata = 32'd20471;
			45066: outdata = 32'd20470;
			45067: outdata = 32'd20469;
			45068: outdata = 32'd20468;
			45069: outdata = 32'd20467;
			45070: outdata = 32'd20466;
			45071: outdata = 32'd20465;
			45072: outdata = 32'd20464;
			45073: outdata = 32'd20463;
			45074: outdata = 32'd20462;
			45075: outdata = 32'd20461;
			45076: outdata = 32'd20460;
			45077: outdata = 32'd20459;
			45078: outdata = 32'd20458;
			45079: outdata = 32'd20457;
			45080: outdata = 32'd20456;
			45081: outdata = 32'd20455;
			45082: outdata = 32'd20454;
			45083: outdata = 32'd20453;
			45084: outdata = 32'd20452;
			45085: outdata = 32'd20451;
			45086: outdata = 32'd20450;
			45087: outdata = 32'd20449;
			45088: outdata = 32'd20448;
			45089: outdata = 32'd20447;
			45090: outdata = 32'd20446;
			45091: outdata = 32'd20445;
			45092: outdata = 32'd20444;
			45093: outdata = 32'd20443;
			45094: outdata = 32'd20442;
			45095: outdata = 32'd20441;
			45096: outdata = 32'd20440;
			45097: outdata = 32'd20439;
			45098: outdata = 32'd20438;
			45099: outdata = 32'd20437;
			45100: outdata = 32'd20436;
			45101: outdata = 32'd20435;
			45102: outdata = 32'd20434;
			45103: outdata = 32'd20433;
			45104: outdata = 32'd20432;
			45105: outdata = 32'd20431;
			45106: outdata = 32'd20430;
			45107: outdata = 32'd20429;
			45108: outdata = 32'd20428;
			45109: outdata = 32'd20427;
			45110: outdata = 32'd20426;
			45111: outdata = 32'd20425;
			45112: outdata = 32'd20424;
			45113: outdata = 32'd20423;
			45114: outdata = 32'd20422;
			45115: outdata = 32'd20421;
			45116: outdata = 32'd20420;
			45117: outdata = 32'd20419;
			45118: outdata = 32'd20418;
			45119: outdata = 32'd20417;
			45120: outdata = 32'd20416;
			45121: outdata = 32'd20415;
			45122: outdata = 32'd20414;
			45123: outdata = 32'd20413;
			45124: outdata = 32'd20412;
			45125: outdata = 32'd20411;
			45126: outdata = 32'd20410;
			45127: outdata = 32'd20409;
			45128: outdata = 32'd20408;
			45129: outdata = 32'd20407;
			45130: outdata = 32'd20406;
			45131: outdata = 32'd20405;
			45132: outdata = 32'd20404;
			45133: outdata = 32'd20403;
			45134: outdata = 32'd20402;
			45135: outdata = 32'd20401;
			45136: outdata = 32'd20400;
			45137: outdata = 32'd20399;
			45138: outdata = 32'd20398;
			45139: outdata = 32'd20397;
			45140: outdata = 32'd20396;
			45141: outdata = 32'd20395;
			45142: outdata = 32'd20394;
			45143: outdata = 32'd20393;
			45144: outdata = 32'd20392;
			45145: outdata = 32'd20391;
			45146: outdata = 32'd20390;
			45147: outdata = 32'd20389;
			45148: outdata = 32'd20388;
			45149: outdata = 32'd20387;
			45150: outdata = 32'd20386;
			45151: outdata = 32'd20385;
			45152: outdata = 32'd20384;
			45153: outdata = 32'd20383;
			45154: outdata = 32'd20382;
			45155: outdata = 32'd20381;
			45156: outdata = 32'd20380;
			45157: outdata = 32'd20379;
			45158: outdata = 32'd20378;
			45159: outdata = 32'd20377;
			45160: outdata = 32'd20376;
			45161: outdata = 32'd20375;
			45162: outdata = 32'd20374;
			45163: outdata = 32'd20373;
			45164: outdata = 32'd20372;
			45165: outdata = 32'd20371;
			45166: outdata = 32'd20370;
			45167: outdata = 32'd20369;
			45168: outdata = 32'd20368;
			45169: outdata = 32'd20367;
			45170: outdata = 32'd20366;
			45171: outdata = 32'd20365;
			45172: outdata = 32'd20364;
			45173: outdata = 32'd20363;
			45174: outdata = 32'd20362;
			45175: outdata = 32'd20361;
			45176: outdata = 32'd20360;
			45177: outdata = 32'd20359;
			45178: outdata = 32'd20358;
			45179: outdata = 32'd20357;
			45180: outdata = 32'd20356;
			45181: outdata = 32'd20355;
			45182: outdata = 32'd20354;
			45183: outdata = 32'd20353;
			45184: outdata = 32'd20352;
			45185: outdata = 32'd20351;
			45186: outdata = 32'd20350;
			45187: outdata = 32'd20349;
			45188: outdata = 32'd20348;
			45189: outdata = 32'd20347;
			45190: outdata = 32'd20346;
			45191: outdata = 32'd20345;
			45192: outdata = 32'd20344;
			45193: outdata = 32'd20343;
			45194: outdata = 32'd20342;
			45195: outdata = 32'd20341;
			45196: outdata = 32'd20340;
			45197: outdata = 32'd20339;
			45198: outdata = 32'd20338;
			45199: outdata = 32'd20337;
			45200: outdata = 32'd20336;
			45201: outdata = 32'd20335;
			45202: outdata = 32'd20334;
			45203: outdata = 32'd20333;
			45204: outdata = 32'd20332;
			45205: outdata = 32'd20331;
			45206: outdata = 32'd20330;
			45207: outdata = 32'd20329;
			45208: outdata = 32'd20328;
			45209: outdata = 32'd20327;
			45210: outdata = 32'd20326;
			45211: outdata = 32'd20325;
			45212: outdata = 32'd20324;
			45213: outdata = 32'd20323;
			45214: outdata = 32'd20322;
			45215: outdata = 32'd20321;
			45216: outdata = 32'd20320;
			45217: outdata = 32'd20319;
			45218: outdata = 32'd20318;
			45219: outdata = 32'd20317;
			45220: outdata = 32'd20316;
			45221: outdata = 32'd20315;
			45222: outdata = 32'd20314;
			45223: outdata = 32'd20313;
			45224: outdata = 32'd20312;
			45225: outdata = 32'd20311;
			45226: outdata = 32'd20310;
			45227: outdata = 32'd20309;
			45228: outdata = 32'd20308;
			45229: outdata = 32'd20307;
			45230: outdata = 32'd20306;
			45231: outdata = 32'd20305;
			45232: outdata = 32'd20304;
			45233: outdata = 32'd20303;
			45234: outdata = 32'd20302;
			45235: outdata = 32'd20301;
			45236: outdata = 32'd20300;
			45237: outdata = 32'd20299;
			45238: outdata = 32'd20298;
			45239: outdata = 32'd20297;
			45240: outdata = 32'd20296;
			45241: outdata = 32'd20295;
			45242: outdata = 32'd20294;
			45243: outdata = 32'd20293;
			45244: outdata = 32'd20292;
			45245: outdata = 32'd20291;
			45246: outdata = 32'd20290;
			45247: outdata = 32'd20289;
			45248: outdata = 32'd20288;
			45249: outdata = 32'd20287;
			45250: outdata = 32'd20286;
			45251: outdata = 32'd20285;
			45252: outdata = 32'd20284;
			45253: outdata = 32'd20283;
			45254: outdata = 32'd20282;
			45255: outdata = 32'd20281;
			45256: outdata = 32'd20280;
			45257: outdata = 32'd20279;
			45258: outdata = 32'd20278;
			45259: outdata = 32'd20277;
			45260: outdata = 32'd20276;
			45261: outdata = 32'd20275;
			45262: outdata = 32'd20274;
			45263: outdata = 32'd20273;
			45264: outdata = 32'd20272;
			45265: outdata = 32'd20271;
			45266: outdata = 32'd20270;
			45267: outdata = 32'd20269;
			45268: outdata = 32'd20268;
			45269: outdata = 32'd20267;
			45270: outdata = 32'd20266;
			45271: outdata = 32'd20265;
			45272: outdata = 32'd20264;
			45273: outdata = 32'd20263;
			45274: outdata = 32'd20262;
			45275: outdata = 32'd20261;
			45276: outdata = 32'd20260;
			45277: outdata = 32'd20259;
			45278: outdata = 32'd20258;
			45279: outdata = 32'd20257;
			45280: outdata = 32'd20256;
			45281: outdata = 32'd20255;
			45282: outdata = 32'd20254;
			45283: outdata = 32'd20253;
			45284: outdata = 32'd20252;
			45285: outdata = 32'd20251;
			45286: outdata = 32'd20250;
			45287: outdata = 32'd20249;
			45288: outdata = 32'd20248;
			45289: outdata = 32'd20247;
			45290: outdata = 32'd20246;
			45291: outdata = 32'd20245;
			45292: outdata = 32'd20244;
			45293: outdata = 32'd20243;
			45294: outdata = 32'd20242;
			45295: outdata = 32'd20241;
			45296: outdata = 32'd20240;
			45297: outdata = 32'd20239;
			45298: outdata = 32'd20238;
			45299: outdata = 32'd20237;
			45300: outdata = 32'd20236;
			45301: outdata = 32'd20235;
			45302: outdata = 32'd20234;
			45303: outdata = 32'd20233;
			45304: outdata = 32'd20232;
			45305: outdata = 32'd20231;
			45306: outdata = 32'd20230;
			45307: outdata = 32'd20229;
			45308: outdata = 32'd20228;
			45309: outdata = 32'd20227;
			45310: outdata = 32'd20226;
			45311: outdata = 32'd20225;
			45312: outdata = 32'd20224;
			45313: outdata = 32'd20223;
			45314: outdata = 32'd20222;
			45315: outdata = 32'd20221;
			45316: outdata = 32'd20220;
			45317: outdata = 32'd20219;
			45318: outdata = 32'd20218;
			45319: outdata = 32'd20217;
			45320: outdata = 32'd20216;
			45321: outdata = 32'd20215;
			45322: outdata = 32'd20214;
			45323: outdata = 32'd20213;
			45324: outdata = 32'd20212;
			45325: outdata = 32'd20211;
			45326: outdata = 32'd20210;
			45327: outdata = 32'd20209;
			45328: outdata = 32'd20208;
			45329: outdata = 32'd20207;
			45330: outdata = 32'd20206;
			45331: outdata = 32'd20205;
			45332: outdata = 32'd20204;
			45333: outdata = 32'd20203;
			45334: outdata = 32'd20202;
			45335: outdata = 32'd20201;
			45336: outdata = 32'd20200;
			45337: outdata = 32'd20199;
			45338: outdata = 32'd20198;
			45339: outdata = 32'd20197;
			45340: outdata = 32'd20196;
			45341: outdata = 32'd20195;
			45342: outdata = 32'd20194;
			45343: outdata = 32'd20193;
			45344: outdata = 32'd20192;
			45345: outdata = 32'd20191;
			45346: outdata = 32'd20190;
			45347: outdata = 32'd20189;
			45348: outdata = 32'd20188;
			45349: outdata = 32'd20187;
			45350: outdata = 32'd20186;
			45351: outdata = 32'd20185;
			45352: outdata = 32'd20184;
			45353: outdata = 32'd20183;
			45354: outdata = 32'd20182;
			45355: outdata = 32'd20181;
			45356: outdata = 32'd20180;
			45357: outdata = 32'd20179;
			45358: outdata = 32'd20178;
			45359: outdata = 32'd20177;
			45360: outdata = 32'd20176;
			45361: outdata = 32'd20175;
			45362: outdata = 32'd20174;
			45363: outdata = 32'd20173;
			45364: outdata = 32'd20172;
			45365: outdata = 32'd20171;
			45366: outdata = 32'd20170;
			45367: outdata = 32'd20169;
			45368: outdata = 32'd20168;
			45369: outdata = 32'd20167;
			45370: outdata = 32'd20166;
			45371: outdata = 32'd20165;
			45372: outdata = 32'd20164;
			45373: outdata = 32'd20163;
			45374: outdata = 32'd20162;
			45375: outdata = 32'd20161;
			45376: outdata = 32'd20160;
			45377: outdata = 32'd20159;
			45378: outdata = 32'd20158;
			45379: outdata = 32'd20157;
			45380: outdata = 32'd20156;
			45381: outdata = 32'd20155;
			45382: outdata = 32'd20154;
			45383: outdata = 32'd20153;
			45384: outdata = 32'd20152;
			45385: outdata = 32'd20151;
			45386: outdata = 32'd20150;
			45387: outdata = 32'd20149;
			45388: outdata = 32'd20148;
			45389: outdata = 32'd20147;
			45390: outdata = 32'd20146;
			45391: outdata = 32'd20145;
			45392: outdata = 32'd20144;
			45393: outdata = 32'd20143;
			45394: outdata = 32'd20142;
			45395: outdata = 32'd20141;
			45396: outdata = 32'd20140;
			45397: outdata = 32'd20139;
			45398: outdata = 32'd20138;
			45399: outdata = 32'd20137;
			45400: outdata = 32'd20136;
			45401: outdata = 32'd20135;
			45402: outdata = 32'd20134;
			45403: outdata = 32'd20133;
			45404: outdata = 32'd20132;
			45405: outdata = 32'd20131;
			45406: outdata = 32'd20130;
			45407: outdata = 32'd20129;
			45408: outdata = 32'd20128;
			45409: outdata = 32'd20127;
			45410: outdata = 32'd20126;
			45411: outdata = 32'd20125;
			45412: outdata = 32'd20124;
			45413: outdata = 32'd20123;
			45414: outdata = 32'd20122;
			45415: outdata = 32'd20121;
			45416: outdata = 32'd20120;
			45417: outdata = 32'd20119;
			45418: outdata = 32'd20118;
			45419: outdata = 32'd20117;
			45420: outdata = 32'd20116;
			45421: outdata = 32'd20115;
			45422: outdata = 32'd20114;
			45423: outdata = 32'd20113;
			45424: outdata = 32'd20112;
			45425: outdata = 32'd20111;
			45426: outdata = 32'd20110;
			45427: outdata = 32'd20109;
			45428: outdata = 32'd20108;
			45429: outdata = 32'd20107;
			45430: outdata = 32'd20106;
			45431: outdata = 32'd20105;
			45432: outdata = 32'd20104;
			45433: outdata = 32'd20103;
			45434: outdata = 32'd20102;
			45435: outdata = 32'd20101;
			45436: outdata = 32'd20100;
			45437: outdata = 32'd20099;
			45438: outdata = 32'd20098;
			45439: outdata = 32'd20097;
			45440: outdata = 32'd20096;
			45441: outdata = 32'd20095;
			45442: outdata = 32'd20094;
			45443: outdata = 32'd20093;
			45444: outdata = 32'd20092;
			45445: outdata = 32'd20091;
			45446: outdata = 32'd20090;
			45447: outdata = 32'd20089;
			45448: outdata = 32'd20088;
			45449: outdata = 32'd20087;
			45450: outdata = 32'd20086;
			45451: outdata = 32'd20085;
			45452: outdata = 32'd20084;
			45453: outdata = 32'd20083;
			45454: outdata = 32'd20082;
			45455: outdata = 32'd20081;
			45456: outdata = 32'd20080;
			45457: outdata = 32'd20079;
			45458: outdata = 32'd20078;
			45459: outdata = 32'd20077;
			45460: outdata = 32'd20076;
			45461: outdata = 32'd20075;
			45462: outdata = 32'd20074;
			45463: outdata = 32'd20073;
			45464: outdata = 32'd20072;
			45465: outdata = 32'd20071;
			45466: outdata = 32'd20070;
			45467: outdata = 32'd20069;
			45468: outdata = 32'd20068;
			45469: outdata = 32'd20067;
			45470: outdata = 32'd20066;
			45471: outdata = 32'd20065;
			45472: outdata = 32'd20064;
			45473: outdata = 32'd20063;
			45474: outdata = 32'd20062;
			45475: outdata = 32'd20061;
			45476: outdata = 32'd20060;
			45477: outdata = 32'd20059;
			45478: outdata = 32'd20058;
			45479: outdata = 32'd20057;
			45480: outdata = 32'd20056;
			45481: outdata = 32'd20055;
			45482: outdata = 32'd20054;
			45483: outdata = 32'd20053;
			45484: outdata = 32'd20052;
			45485: outdata = 32'd20051;
			45486: outdata = 32'd20050;
			45487: outdata = 32'd20049;
			45488: outdata = 32'd20048;
			45489: outdata = 32'd20047;
			45490: outdata = 32'd20046;
			45491: outdata = 32'd20045;
			45492: outdata = 32'd20044;
			45493: outdata = 32'd20043;
			45494: outdata = 32'd20042;
			45495: outdata = 32'd20041;
			45496: outdata = 32'd20040;
			45497: outdata = 32'd20039;
			45498: outdata = 32'd20038;
			45499: outdata = 32'd20037;
			45500: outdata = 32'd20036;
			45501: outdata = 32'd20035;
			45502: outdata = 32'd20034;
			45503: outdata = 32'd20033;
			45504: outdata = 32'd20032;
			45505: outdata = 32'd20031;
			45506: outdata = 32'd20030;
			45507: outdata = 32'd20029;
			45508: outdata = 32'd20028;
			45509: outdata = 32'd20027;
			45510: outdata = 32'd20026;
			45511: outdata = 32'd20025;
			45512: outdata = 32'd20024;
			45513: outdata = 32'd20023;
			45514: outdata = 32'd20022;
			45515: outdata = 32'd20021;
			45516: outdata = 32'd20020;
			45517: outdata = 32'd20019;
			45518: outdata = 32'd20018;
			45519: outdata = 32'd20017;
			45520: outdata = 32'd20016;
			45521: outdata = 32'd20015;
			45522: outdata = 32'd20014;
			45523: outdata = 32'd20013;
			45524: outdata = 32'd20012;
			45525: outdata = 32'd20011;
			45526: outdata = 32'd20010;
			45527: outdata = 32'd20009;
			45528: outdata = 32'd20008;
			45529: outdata = 32'd20007;
			45530: outdata = 32'd20006;
			45531: outdata = 32'd20005;
			45532: outdata = 32'd20004;
			45533: outdata = 32'd20003;
			45534: outdata = 32'd20002;
			45535: outdata = 32'd20001;
			45536: outdata = 32'd20000;
			45537: outdata = 32'd19999;
			45538: outdata = 32'd19998;
			45539: outdata = 32'd19997;
			45540: outdata = 32'd19996;
			45541: outdata = 32'd19995;
			45542: outdata = 32'd19994;
			45543: outdata = 32'd19993;
			45544: outdata = 32'd19992;
			45545: outdata = 32'd19991;
			45546: outdata = 32'd19990;
			45547: outdata = 32'd19989;
			45548: outdata = 32'd19988;
			45549: outdata = 32'd19987;
			45550: outdata = 32'd19986;
			45551: outdata = 32'd19985;
			45552: outdata = 32'd19984;
			45553: outdata = 32'd19983;
			45554: outdata = 32'd19982;
			45555: outdata = 32'd19981;
			45556: outdata = 32'd19980;
			45557: outdata = 32'd19979;
			45558: outdata = 32'd19978;
			45559: outdata = 32'd19977;
			45560: outdata = 32'd19976;
			45561: outdata = 32'd19975;
			45562: outdata = 32'd19974;
			45563: outdata = 32'd19973;
			45564: outdata = 32'd19972;
			45565: outdata = 32'd19971;
			45566: outdata = 32'd19970;
			45567: outdata = 32'd19969;
			45568: outdata = 32'd19968;
			45569: outdata = 32'd19967;
			45570: outdata = 32'd19966;
			45571: outdata = 32'd19965;
			45572: outdata = 32'd19964;
			45573: outdata = 32'd19963;
			45574: outdata = 32'd19962;
			45575: outdata = 32'd19961;
			45576: outdata = 32'd19960;
			45577: outdata = 32'd19959;
			45578: outdata = 32'd19958;
			45579: outdata = 32'd19957;
			45580: outdata = 32'd19956;
			45581: outdata = 32'd19955;
			45582: outdata = 32'd19954;
			45583: outdata = 32'd19953;
			45584: outdata = 32'd19952;
			45585: outdata = 32'd19951;
			45586: outdata = 32'd19950;
			45587: outdata = 32'd19949;
			45588: outdata = 32'd19948;
			45589: outdata = 32'd19947;
			45590: outdata = 32'd19946;
			45591: outdata = 32'd19945;
			45592: outdata = 32'd19944;
			45593: outdata = 32'd19943;
			45594: outdata = 32'd19942;
			45595: outdata = 32'd19941;
			45596: outdata = 32'd19940;
			45597: outdata = 32'd19939;
			45598: outdata = 32'd19938;
			45599: outdata = 32'd19937;
			45600: outdata = 32'd19936;
			45601: outdata = 32'd19935;
			45602: outdata = 32'd19934;
			45603: outdata = 32'd19933;
			45604: outdata = 32'd19932;
			45605: outdata = 32'd19931;
			45606: outdata = 32'd19930;
			45607: outdata = 32'd19929;
			45608: outdata = 32'd19928;
			45609: outdata = 32'd19927;
			45610: outdata = 32'd19926;
			45611: outdata = 32'd19925;
			45612: outdata = 32'd19924;
			45613: outdata = 32'd19923;
			45614: outdata = 32'd19922;
			45615: outdata = 32'd19921;
			45616: outdata = 32'd19920;
			45617: outdata = 32'd19919;
			45618: outdata = 32'd19918;
			45619: outdata = 32'd19917;
			45620: outdata = 32'd19916;
			45621: outdata = 32'd19915;
			45622: outdata = 32'd19914;
			45623: outdata = 32'd19913;
			45624: outdata = 32'd19912;
			45625: outdata = 32'd19911;
			45626: outdata = 32'd19910;
			45627: outdata = 32'd19909;
			45628: outdata = 32'd19908;
			45629: outdata = 32'd19907;
			45630: outdata = 32'd19906;
			45631: outdata = 32'd19905;
			45632: outdata = 32'd19904;
			45633: outdata = 32'd19903;
			45634: outdata = 32'd19902;
			45635: outdata = 32'd19901;
			45636: outdata = 32'd19900;
			45637: outdata = 32'd19899;
			45638: outdata = 32'd19898;
			45639: outdata = 32'd19897;
			45640: outdata = 32'd19896;
			45641: outdata = 32'd19895;
			45642: outdata = 32'd19894;
			45643: outdata = 32'd19893;
			45644: outdata = 32'd19892;
			45645: outdata = 32'd19891;
			45646: outdata = 32'd19890;
			45647: outdata = 32'd19889;
			45648: outdata = 32'd19888;
			45649: outdata = 32'd19887;
			45650: outdata = 32'd19886;
			45651: outdata = 32'd19885;
			45652: outdata = 32'd19884;
			45653: outdata = 32'd19883;
			45654: outdata = 32'd19882;
			45655: outdata = 32'd19881;
			45656: outdata = 32'd19880;
			45657: outdata = 32'd19879;
			45658: outdata = 32'd19878;
			45659: outdata = 32'd19877;
			45660: outdata = 32'd19876;
			45661: outdata = 32'd19875;
			45662: outdata = 32'd19874;
			45663: outdata = 32'd19873;
			45664: outdata = 32'd19872;
			45665: outdata = 32'd19871;
			45666: outdata = 32'd19870;
			45667: outdata = 32'd19869;
			45668: outdata = 32'd19868;
			45669: outdata = 32'd19867;
			45670: outdata = 32'd19866;
			45671: outdata = 32'd19865;
			45672: outdata = 32'd19864;
			45673: outdata = 32'd19863;
			45674: outdata = 32'd19862;
			45675: outdata = 32'd19861;
			45676: outdata = 32'd19860;
			45677: outdata = 32'd19859;
			45678: outdata = 32'd19858;
			45679: outdata = 32'd19857;
			45680: outdata = 32'd19856;
			45681: outdata = 32'd19855;
			45682: outdata = 32'd19854;
			45683: outdata = 32'd19853;
			45684: outdata = 32'd19852;
			45685: outdata = 32'd19851;
			45686: outdata = 32'd19850;
			45687: outdata = 32'd19849;
			45688: outdata = 32'd19848;
			45689: outdata = 32'd19847;
			45690: outdata = 32'd19846;
			45691: outdata = 32'd19845;
			45692: outdata = 32'd19844;
			45693: outdata = 32'd19843;
			45694: outdata = 32'd19842;
			45695: outdata = 32'd19841;
			45696: outdata = 32'd19840;
			45697: outdata = 32'd19839;
			45698: outdata = 32'd19838;
			45699: outdata = 32'd19837;
			45700: outdata = 32'd19836;
			45701: outdata = 32'd19835;
			45702: outdata = 32'd19834;
			45703: outdata = 32'd19833;
			45704: outdata = 32'd19832;
			45705: outdata = 32'd19831;
			45706: outdata = 32'd19830;
			45707: outdata = 32'd19829;
			45708: outdata = 32'd19828;
			45709: outdata = 32'd19827;
			45710: outdata = 32'd19826;
			45711: outdata = 32'd19825;
			45712: outdata = 32'd19824;
			45713: outdata = 32'd19823;
			45714: outdata = 32'd19822;
			45715: outdata = 32'd19821;
			45716: outdata = 32'd19820;
			45717: outdata = 32'd19819;
			45718: outdata = 32'd19818;
			45719: outdata = 32'd19817;
			45720: outdata = 32'd19816;
			45721: outdata = 32'd19815;
			45722: outdata = 32'd19814;
			45723: outdata = 32'd19813;
			45724: outdata = 32'd19812;
			45725: outdata = 32'd19811;
			45726: outdata = 32'd19810;
			45727: outdata = 32'd19809;
			45728: outdata = 32'd19808;
			45729: outdata = 32'd19807;
			45730: outdata = 32'd19806;
			45731: outdata = 32'd19805;
			45732: outdata = 32'd19804;
			45733: outdata = 32'd19803;
			45734: outdata = 32'd19802;
			45735: outdata = 32'd19801;
			45736: outdata = 32'd19800;
			45737: outdata = 32'd19799;
			45738: outdata = 32'd19798;
			45739: outdata = 32'd19797;
			45740: outdata = 32'd19796;
			45741: outdata = 32'd19795;
			45742: outdata = 32'd19794;
			45743: outdata = 32'd19793;
			45744: outdata = 32'd19792;
			45745: outdata = 32'd19791;
			45746: outdata = 32'd19790;
			45747: outdata = 32'd19789;
			45748: outdata = 32'd19788;
			45749: outdata = 32'd19787;
			45750: outdata = 32'd19786;
			45751: outdata = 32'd19785;
			45752: outdata = 32'd19784;
			45753: outdata = 32'd19783;
			45754: outdata = 32'd19782;
			45755: outdata = 32'd19781;
			45756: outdata = 32'd19780;
			45757: outdata = 32'd19779;
			45758: outdata = 32'd19778;
			45759: outdata = 32'd19777;
			45760: outdata = 32'd19776;
			45761: outdata = 32'd19775;
			45762: outdata = 32'd19774;
			45763: outdata = 32'd19773;
			45764: outdata = 32'd19772;
			45765: outdata = 32'd19771;
			45766: outdata = 32'd19770;
			45767: outdata = 32'd19769;
			45768: outdata = 32'd19768;
			45769: outdata = 32'd19767;
			45770: outdata = 32'd19766;
			45771: outdata = 32'd19765;
			45772: outdata = 32'd19764;
			45773: outdata = 32'd19763;
			45774: outdata = 32'd19762;
			45775: outdata = 32'd19761;
			45776: outdata = 32'd19760;
			45777: outdata = 32'd19759;
			45778: outdata = 32'd19758;
			45779: outdata = 32'd19757;
			45780: outdata = 32'd19756;
			45781: outdata = 32'd19755;
			45782: outdata = 32'd19754;
			45783: outdata = 32'd19753;
			45784: outdata = 32'd19752;
			45785: outdata = 32'd19751;
			45786: outdata = 32'd19750;
			45787: outdata = 32'd19749;
			45788: outdata = 32'd19748;
			45789: outdata = 32'd19747;
			45790: outdata = 32'd19746;
			45791: outdata = 32'd19745;
			45792: outdata = 32'd19744;
			45793: outdata = 32'd19743;
			45794: outdata = 32'd19742;
			45795: outdata = 32'd19741;
			45796: outdata = 32'd19740;
			45797: outdata = 32'd19739;
			45798: outdata = 32'd19738;
			45799: outdata = 32'd19737;
			45800: outdata = 32'd19736;
			45801: outdata = 32'd19735;
			45802: outdata = 32'd19734;
			45803: outdata = 32'd19733;
			45804: outdata = 32'd19732;
			45805: outdata = 32'd19731;
			45806: outdata = 32'd19730;
			45807: outdata = 32'd19729;
			45808: outdata = 32'd19728;
			45809: outdata = 32'd19727;
			45810: outdata = 32'd19726;
			45811: outdata = 32'd19725;
			45812: outdata = 32'd19724;
			45813: outdata = 32'd19723;
			45814: outdata = 32'd19722;
			45815: outdata = 32'd19721;
			45816: outdata = 32'd19720;
			45817: outdata = 32'd19719;
			45818: outdata = 32'd19718;
			45819: outdata = 32'd19717;
			45820: outdata = 32'd19716;
			45821: outdata = 32'd19715;
			45822: outdata = 32'd19714;
			45823: outdata = 32'd19713;
			45824: outdata = 32'd19712;
			45825: outdata = 32'd19711;
			45826: outdata = 32'd19710;
			45827: outdata = 32'd19709;
			45828: outdata = 32'd19708;
			45829: outdata = 32'd19707;
			45830: outdata = 32'd19706;
			45831: outdata = 32'd19705;
			45832: outdata = 32'd19704;
			45833: outdata = 32'd19703;
			45834: outdata = 32'd19702;
			45835: outdata = 32'd19701;
			45836: outdata = 32'd19700;
			45837: outdata = 32'd19699;
			45838: outdata = 32'd19698;
			45839: outdata = 32'd19697;
			45840: outdata = 32'd19696;
			45841: outdata = 32'd19695;
			45842: outdata = 32'd19694;
			45843: outdata = 32'd19693;
			45844: outdata = 32'd19692;
			45845: outdata = 32'd19691;
			45846: outdata = 32'd19690;
			45847: outdata = 32'd19689;
			45848: outdata = 32'd19688;
			45849: outdata = 32'd19687;
			45850: outdata = 32'd19686;
			45851: outdata = 32'd19685;
			45852: outdata = 32'd19684;
			45853: outdata = 32'd19683;
			45854: outdata = 32'd19682;
			45855: outdata = 32'd19681;
			45856: outdata = 32'd19680;
			45857: outdata = 32'd19679;
			45858: outdata = 32'd19678;
			45859: outdata = 32'd19677;
			45860: outdata = 32'd19676;
			45861: outdata = 32'd19675;
			45862: outdata = 32'd19674;
			45863: outdata = 32'd19673;
			45864: outdata = 32'd19672;
			45865: outdata = 32'd19671;
			45866: outdata = 32'd19670;
			45867: outdata = 32'd19669;
			45868: outdata = 32'd19668;
			45869: outdata = 32'd19667;
			45870: outdata = 32'd19666;
			45871: outdata = 32'd19665;
			45872: outdata = 32'd19664;
			45873: outdata = 32'd19663;
			45874: outdata = 32'd19662;
			45875: outdata = 32'd19661;
			45876: outdata = 32'd19660;
			45877: outdata = 32'd19659;
			45878: outdata = 32'd19658;
			45879: outdata = 32'd19657;
			45880: outdata = 32'd19656;
			45881: outdata = 32'd19655;
			45882: outdata = 32'd19654;
			45883: outdata = 32'd19653;
			45884: outdata = 32'd19652;
			45885: outdata = 32'd19651;
			45886: outdata = 32'd19650;
			45887: outdata = 32'd19649;
			45888: outdata = 32'd19648;
			45889: outdata = 32'd19647;
			45890: outdata = 32'd19646;
			45891: outdata = 32'd19645;
			45892: outdata = 32'd19644;
			45893: outdata = 32'd19643;
			45894: outdata = 32'd19642;
			45895: outdata = 32'd19641;
			45896: outdata = 32'd19640;
			45897: outdata = 32'd19639;
			45898: outdata = 32'd19638;
			45899: outdata = 32'd19637;
			45900: outdata = 32'd19636;
			45901: outdata = 32'd19635;
			45902: outdata = 32'd19634;
			45903: outdata = 32'd19633;
			45904: outdata = 32'd19632;
			45905: outdata = 32'd19631;
			45906: outdata = 32'd19630;
			45907: outdata = 32'd19629;
			45908: outdata = 32'd19628;
			45909: outdata = 32'd19627;
			45910: outdata = 32'd19626;
			45911: outdata = 32'd19625;
			45912: outdata = 32'd19624;
			45913: outdata = 32'd19623;
			45914: outdata = 32'd19622;
			45915: outdata = 32'd19621;
			45916: outdata = 32'd19620;
			45917: outdata = 32'd19619;
			45918: outdata = 32'd19618;
			45919: outdata = 32'd19617;
			45920: outdata = 32'd19616;
			45921: outdata = 32'd19615;
			45922: outdata = 32'd19614;
			45923: outdata = 32'd19613;
			45924: outdata = 32'd19612;
			45925: outdata = 32'd19611;
			45926: outdata = 32'd19610;
			45927: outdata = 32'd19609;
			45928: outdata = 32'd19608;
			45929: outdata = 32'd19607;
			45930: outdata = 32'd19606;
			45931: outdata = 32'd19605;
			45932: outdata = 32'd19604;
			45933: outdata = 32'd19603;
			45934: outdata = 32'd19602;
			45935: outdata = 32'd19601;
			45936: outdata = 32'd19600;
			45937: outdata = 32'd19599;
			45938: outdata = 32'd19598;
			45939: outdata = 32'd19597;
			45940: outdata = 32'd19596;
			45941: outdata = 32'd19595;
			45942: outdata = 32'd19594;
			45943: outdata = 32'd19593;
			45944: outdata = 32'd19592;
			45945: outdata = 32'd19591;
			45946: outdata = 32'd19590;
			45947: outdata = 32'd19589;
			45948: outdata = 32'd19588;
			45949: outdata = 32'd19587;
			45950: outdata = 32'd19586;
			45951: outdata = 32'd19585;
			45952: outdata = 32'd19584;
			45953: outdata = 32'd19583;
			45954: outdata = 32'd19582;
			45955: outdata = 32'd19581;
			45956: outdata = 32'd19580;
			45957: outdata = 32'd19579;
			45958: outdata = 32'd19578;
			45959: outdata = 32'd19577;
			45960: outdata = 32'd19576;
			45961: outdata = 32'd19575;
			45962: outdata = 32'd19574;
			45963: outdata = 32'd19573;
			45964: outdata = 32'd19572;
			45965: outdata = 32'd19571;
			45966: outdata = 32'd19570;
			45967: outdata = 32'd19569;
			45968: outdata = 32'd19568;
			45969: outdata = 32'd19567;
			45970: outdata = 32'd19566;
			45971: outdata = 32'd19565;
			45972: outdata = 32'd19564;
			45973: outdata = 32'd19563;
			45974: outdata = 32'd19562;
			45975: outdata = 32'd19561;
			45976: outdata = 32'd19560;
			45977: outdata = 32'd19559;
			45978: outdata = 32'd19558;
			45979: outdata = 32'd19557;
			45980: outdata = 32'd19556;
			45981: outdata = 32'd19555;
			45982: outdata = 32'd19554;
			45983: outdata = 32'd19553;
			45984: outdata = 32'd19552;
			45985: outdata = 32'd19551;
			45986: outdata = 32'd19550;
			45987: outdata = 32'd19549;
			45988: outdata = 32'd19548;
			45989: outdata = 32'd19547;
			45990: outdata = 32'd19546;
			45991: outdata = 32'd19545;
			45992: outdata = 32'd19544;
			45993: outdata = 32'd19543;
			45994: outdata = 32'd19542;
			45995: outdata = 32'd19541;
			45996: outdata = 32'd19540;
			45997: outdata = 32'd19539;
			45998: outdata = 32'd19538;
			45999: outdata = 32'd19537;
			46000: outdata = 32'd19536;
			46001: outdata = 32'd19535;
			46002: outdata = 32'd19534;
			46003: outdata = 32'd19533;
			46004: outdata = 32'd19532;
			46005: outdata = 32'd19531;
			46006: outdata = 32'd19530;
			46007: outdata = 32'd19529;
			46008: outdata = 32'd19528;
			46009: outdata = 32'd19527;
			46010: outdata = 32'd19526;
			46011: outdata = 32'd19525;
			46012: outdata = 32'd19524;
			46013: outdata = 32'd19523;
			46014: outdata = 32'd19522;
			46015: outdata = 32'd19521;
			46016: outdata = 32'd19520;
			46017: outdata = 32'd19519;
			46018: outdata = 32'd19518;
			46019: outdata = 32'd19517;
			46020: outdata = 32'd19516;
			46021: outdata = 32'd19515;
			46022: outdata = 32'd19514;
			46023: outdata = 32'd19513;
			46024: outdata = 32'd19512;
			46025: outdata = 32'd19511;
			46026: outdata = 32'd19510;
			46027: outdata = 32'd19509;
			46028: outdata = 32'd19508;
			46029: outdata = 32'd19507;
			46030: outdata = 32'd19506;
			46031: outdata = 32'd19505;
			46032: outdata = 32'd19504;
			46033: outdata = 32'd19503;
			46034: outdata = 32'd19502;
			46035: outdata = 32'd19501;
			46036: outdata = 32'd19500;
			46037: outdata = 32'd19499;
			46038: outdata = 32'd19498;
			46039: outdata = 32'd19497;
			46040: outdata = 32'd19496;
			46041: outdata = 32'd19495;
			46042: outdata = 32'd19494;
			46043: outdata = 32'd19493;
			46044: outdata = 32'd19492;
			46045: outdata = 32'd19491;
			46046: outdata = 32'd19490;
			46047: outdata = 32'd19489;
			46048: outdata = 32'd19488;
			46049: outdata = 32'd19487;
			46050: outdata = 32'd19486;
			46051: outdata = 32'd19485;
			46052: outdata = 32'd19484;
			46053: outdata = 32'd19483;
			46054: outdata = 32'd19482;
			46055: outdata = 32'd19481;
			46056: outdata = 32'd19480;
			46057: outdata = 32'd19479;
			46058: outdata = 32'd19478;
			46059: outdata = 32'd19477;
			46060: outdata = 32'd19476;
			46061: outdata = 32'd19475;
			46062: outdata = 32'd19474;
			46063: outdata = 32'd19473;
			46064: outdata = 32'd19472;
			46065: outdata = 32'd19471;
			46066: outdata = 32'd19470;
			46067: outdata = 32'd19469;
			46068: outdata = 32'd19468;
			46069: outdata = 32'd19467;
			46070: outdata = 32'd19466;
			46071: outdata = 32'd19465;
			46072: outdata = 32'd19464;
			46073: outdata = 32'd19463;
			46074: outdata = 32'd19462;
			46075: outdata = 32'd19461;
			46076: outdata = 32'd19460;
			46077: outdata = 32'd19459;
			46078: outdata = 32'd19458;
			46079: outdata = 32'd19457;
			46080: outdata = 32'd19456;
			46081: outdata = 32'd19455;
			46082: outdata = 32'd19454;
			46083: outdata = 32'd19453;
			46084: outdata = 32'd19452;
			46085: outdata = 32'd19451;
			46086: outdata = 32'd19450;
			46087: outdata = 32'd19449;
			46088: outdata = 32'd19448;
			46089: outdata = 32'd19447;
			46090: outdata = 32'd19446;
			46091: outdata = 32'd19445;
			46092: outdata = 32'd19444;
			46093: outdata = 32'd19443;
			46094: outdata = 32'd19442;
			46095: outdata = 32'd19441;
			46096: outdata = 32'd19440;
			46097: outdata = 32'd19439;
			46098: outdata = 32'd19438;
			46099: outdata = 32'd19437;
			46100: outdata = 32'd19436;
			46101: outdata = 32'd19435;
			46102: outdata = 32'd19434;
			46103: outdata = 32'd19433;
			46104: outdata = 32'd19432;
			46105: outdata = 32'd19431;
			46106: outdata = 32'd19430;
			46107: outdata = 32'd19429;
			46108: outdata = 32'd19428;
			46109: outdata = 32'd19427;
			46110: outdata = 32'd19426;
			46111: outdata = 32'd19425;
			46112: outdata = 32'd19424;
			46113: outdata = 32'd19423;
			46114: outdata = 32'd19422;
			46115: outdata = 32'd19421;
			46116: outdata = 32'd19420;
			46117: outdata = 32'd19419;
			46118: outdata = 32'd19418;
			46119: outdata = 32'd19417;
			46120: outdata = 32'd19416;
			46121: outdata = 32'd19415;
			46122: outdata = 32'd19414;
			46123: outdata = 32'd19413;
			46124: outdata = 32'd19412;
			46125: outdata = 32'd19411;
			46126: outdata = 32'd19410;
			46127: outdata = 32'd19409;
			46128: outdata = 32'd19408;
			46129: outdata = 32'd19407;
			46130: outdata = 32'd19406;
			46131: outdata = 32'd19405;
			46132: outdata = 32'd19404;
			46133: outdata = 32'd19403;
			46134: outdata = 32'd19402;
			46135: outdata = 32'd19401;
			46136: outdata = 32'd19400;
			46137: outdata = 32'd19399;
			46138: outdata = 32'd19398;
			46139: outdata = 32'd19397;
			46140: outdata = 32'd19396;
			46141: outdata = 32'd19395;
			46142: outdata = 32'd19394;
			46143: outdata = 32'd19393;
			46144: outdata = 32'd19392;
			46145: outdata = 32'd19391;
			46146: outdata = 32'd19390;
			46147: outdata = 32'd19389;
			46148: outdata = 32'd19388;
			46149: outdata = 32'd19387;
			46150: outdata = 32'd19386;
			46151: outdata = 32'd19385;
			46152: outdata = 32'd19384;
			46153: outdata = 32'd19383;
			46154: outdata = 32'd19382;
			46155: outdata = 32'd19381;
			46156: outdata = 32'd19380;
			46157: outdata = 32'd19379;
			46158: outdata = 32'd19378;
			46159: outdata = 32'd19377;
			46160: outdata = 32'd19376;
			46161: outdata = 32'd19375;
			46162: outdata = 32'd19374;
			46163: outdata = 32'd19373;
			46164: outdata = 32'd19372;
			46165: outdata = 32'd19371;
			46166: outdata = 32'd19370;
			46167: outdata = 32'd19369;
			46168: outdata = 32'd19368;
			46169: outdata = 32'd19367;
			46170: outdata = 32'd19366;
			46171: outdata = 32'd19365;
			46172: outdata = 32'd19364;
			46173: outdata = 32'd19363;
			46174: outdata = 32'd19362;
			46175: outdata = 32'd19361;
			46176: outdata = 32'd19360;
			46177: outdata = 32'd19359;
			46178: outdata = 32'd19358;
			46179: outdata = 32'd19357;
			46180: outdata = 32'd19356;
			46181: outdata = 32'd19355;
			46182: outdata = 32'd19354;
			46183: outdata = 32'd19353;
			46184: outdata = 32'd19352;
			46185: outdata = 32'd19351;
			46186: outdata = 32'd19350;
			46187: outdata = 32'd19349;
			46188: outdata = 32'd19348;
			46189: outdata = 32'd19347;
			46190: outdata = 32'd19346;
			46191: outdata = 32'd19345;
			46192: outdata = 32'd19344;
			46193: outdata = 32'd19343;
			46194: outdata = 32'd19342;
			46195: outdata = 32'd19341;
			46196: outdata = 32'd19340;
			46197: outdata = 32'd19339;
			46198: outdata = 32'd19338;
			46199: outdata = 32'd19337;
			46200: outdata = 32'd19336;
			46201: outdata = 32'd19335;
			46202: outdata = 32'd19334;
			46203: outdata = 32'd19333;
			46204: outdata = 32'd19332;
			46205: outdata = 32'd19331;
			46206: outdata = 32'd19330;
			46207: outdata = 32'd19329;
			46208: outdata = 32'd19328;
			46209: outdata = 32'd19327;
			46210: outdata = 32'd19326;
			46211: outdata = 32'd19325;
			46212: outdata = 32'd19324;
			46213: outdata = 32'd19323;
			46214: outdata = 32'd19322;
			46215: outdata = 32'd19321;
			46216: outdata = 32'd19320;
			46217: outdata = 32'd19319;
			46218: outdata = 32'd19318;
			46219: outdata = 32'd19317;
			46220: outdata = 32'd19316;
			46221: outdata = 32'd19315;
			46222: outdata = 32'd19314;
			46223: outdata = 32'd19313;
			46224: outdata = 32'd19312;
			46225: outdata = 32'd19311;
			46226: outdata = 32'd19310;
			46227: outdata = 32'd19309;
			46228: outdata = 32'd19308;
			46229: outdata = 32'd19307;
			46230: outdata = 32'd19306;
			46231: outdata = 32'd19305;
			46232: outdata = 32'd19304;
			46233: outdata = 32'd19303;
			46234: outdata = 32'd19302;
			46235: outdata = 32'd19301;
			46236: outdata = 32'd19300;
			46237: outdata = 32'd19299;
			46238: outdata = 32'd19298;
			46239: outdata = 32'd19297;
			46240: outdata = 32'd19296;
			46241: outdata = 32'd19295;
			46242: outdata = 32'd19294;
			46243: outdata = 32'd19293;
			46244: outdata = 32'd19292;
			46245: outdata = 32'd19291;
			46246: outdata = 32'd19290;
			46247: outdata = 32'd19289;
			46248: outdata = 32'd19288;
			46249: outdata = 32'd19287;
			46250: outdata = 32'd19286;
			46251: outdata = 32'd19285;
			46252: outdata = 32'd19284;
			46253: outdata = 32'd19283;
			46254: outdata = 32'd19282;
			46255: outdata = 32'd19281;
			46256: outdata = 32'd19280;
			46257: outdata = 32'd19279;
			46258: outdata = 32'd19278;
			46259: outdata = 32'd19277;
			46260: outdata = 32'd19276;
			46261: outdata = 32'd19275;
			46262: outdata = 32'd19274;
			46263: outdata = 32'd19273;
			46264: outdata = 32'd19272;
			46265: outdata = 32'd19271;
			46266: outdata = 32'd19270;
			46267: outdata = 32'd19269;
			46268: outdata = 32'd19268;
			46269: outdata = 32'd19267;
			46270: outdata = 32'd19266;
			46271: outdata = 32'd19265;
			46272: outdata = 32'd19264;
			46273: outdata = 32'd19263;
			46274: outdata = 32'd19262;
			46275: outdata = 32'd19261;
			46276: outdata = 32'd19260;
			46277: outdata = 32'd19259;
			46278: outdata = 32'd19258;
			46279: outdata = 32'd19257;
			46280: outdata = 32'd19256;
			46281: outdata = 32'd19255;
			46282: outdata = 32'd19254;
			46283: outdata = 32'd19253;
			46284: outdata = 32'd19252;
			46285: outdata = 32'd19251;
			46286: outdata = 32'd19250;
			46287: outdata = 32'd19249;
			46288: outdata = 32'd19248;
			46289: outdata = 32'd19247;
			46290: outdata = 32'd19246;
			46291: outdata = 32'd19245;
			46292: outdata = 32'd19244;
			46293: outdata = 32'd19243;
			46294: outdata = 32'd19242;
			46295: outdata = 32'd19241;
			46296: outdata = 32'd19240;
			46297: outdata = 32'd19239;
			46298: outdata = 32'd19238;
			46299: outdata = 32'd19237;
			46300: outdata = 32'd19236;
			46301: outdata = 32'd19235;
			46302: outdata = 32'd19234;
			46303: outdata = 32'd19233;
			46304: outdata = 32'd19232;
			46305: outdata = 32'd19231;
			46306: outdata = 32'd19230;
			46307: outdata = 32'd19229;
			46308: outdata = 32'd19228;
			46309: outdata = 32'd19227;
			46310: outdata = 32'd19226;
			46311: outdata = 32'd19225;
			46312: outdata = 32'd19224;
			46313: outdata = 32'd19223;
			46314: outdata = 32'd19222;
			46315: outdata = 32'd19221;
			46316: outdata = 32'd19220;
			46317: outdata = 32'd19219;
			46318: outdata = 32'd19218;
			46319: outdata = 32'd19217;
			46320: outdata = 32'd19216;
			46321: outdata = 32'd19215;
			46322: outdata = 32'd19214;
			46323: outdata = 32'd19213;
			46324: outdata = 32'd19212;
			46325: outdata = 32'd19211;
			46326: outdata = 32'd19210;
			46327: outdata = 32'd19209;
			46328: outdata = 32'd19208;
			46329: outdata = 32'd19207;
			46330: outdata = 32'd19206;
			46331: outdata = 32'd19205;
			46332: outdata = 32'd19204;
			46333: outdata = 32'd19203;
			46334: outdata = 32'd19202;
			46335: outdata = 32'd19201;
			46336: outdata = 32'd19200;
			46337: outdata = 32'd19199;
			46338: outdata = 32'd19198;
			46339: outdata = 32'd19197;
			46340: outdata = 32'd19196;
			46341: outdata = 32'd19195;
			46342: outdata = 32'd19194;
			46343: outdata = 32'd19193;
			46344: outdata = 32'd19192;
			46345: outdata = 32'd19191;
			46346: outdata = 32'd19190;
			46347: outdata = 32'd19189;
			46348: outdata = 32'd19188;
			46349: outdata = 32'd19187;
			46350: outdata = 32'd19186;
			46351: outdata = 32'd19185;
			46352: outdata = 32'd19184;
			46353: outdata = 32'd19183;
			46354: outdata = 32'd19182;
			46355: outdata = 32'd19181;
			46356: outdata = 32'd19180;
			46357: outdata = 32'd19179;
			46358: outdata = 32'd19178;
			46359: outdata = 32'd19177;
			46360: outdata = 32'd19176;
			46361: outdata = 32'd19175;
			46362: outdata = 32'd19174;
			46363: outdata = 32'd19173;
			46364: outdata = 32'd19172;
			46365: outdata = 32'd19171;
			46366: outdata = 32'd19170;
			46367: outdata = 32'd19169;
			46368: outdata = 32'd19168;
			46369: outdata = 32'd19167;
			46370: outdata = 32'd19166;
			46371: outdata = 32'd19165;
			46372: outdata = 32'd19164;
			46373: outdata = 32'd19163;
			46374: outdata = 32'd19162;
			46375: outdata = 32'd19161;
			46376: outdata = 32'd19160;
			46377: outdata = 32'd19159;
			46378: outdata = 32'd19158;
			46379: outdata = 32'd19157;
			46380: outdata = 32'd19156;
			46381: outdata = 32'd19155;
			46382: outdata = 32'd19154;
			46383: outdata = 32'd19153;
			46384: outdata = 32'd19152;
			46385: outdata = 32'd19151;
			46386: outdata = 32'd19150;
			46387: outdata = 32'd19149;
			46388: outdata = 32'd19148;
			46389: outdata = 32'd19147;
			46390: outdata = 32'd19146;
			46391: outdata = 32'd19145;
			46392: outdata = 32'd19144;
			46393: outdata = 32'd19143;
			46394: outdata = 32'd19142;
			46395: outdata = 32'd19141;
			46396: outdata = 32'd19140;
			46397: outdata = 32'd19139;
			46398: outdata = 32'd19138;
			46399: outdata = 32'd19137;
			46400: outdata = 32'd19136;
			46401: outdata = 32'd19135;
			46402: outdata = 32'd19134;
			46403: outdata = 32'd19133;
			46404: outdata = 32'd19132;
			46405: outdata = 32'd19131;
			46406: outdata = 32'd19130;
			46407: outdata = 32'd19129;
			46408: outdata = 32'd19128;
			46409: outdata = 32'd19127;
			46410: outdata = 32'd19126;
			46411: outdata = 32'd19125;
			46412: outdata = 32'd19124;
			46413: outdata = 32'd19123;
			46414: outdata = 32'd19122;
			46415: outdata = 32'd19121;
			46416: outdata = 32'd19120;
			46417: outdata = 32'd19119;
			46418: outdata = 32'd19118;
			46419: outdata = 32'd19117;
			46420: outdata = 32'd19116;
			46421: outdata = 32'd19115;
			46422: outdata = 32'd19114;
			46423: outdata = 32'd19113;
			46424: outdata = 32'd19112;
			46425: outdata = 32'd19111;
			46426: outdata = 32'd19110;
			46427: outdata = 32'd19109;
			46428: outdata = 32'd19108;
			46429: outdata = 32'd19107;
			46430: outdata = 32'd19106;
			46431: outdata = 32'd19105;
			46432: outdata = 32'd19104;
			46433: outdata = 32'd19103;
			46434: outdata = 32'd19102;
			46435: outdata = 32'd19101;
			46436: outdata = 32'd19100;
			46437: outdata = 32'd19099;
			46438: outdata = 32'd19098;
			46439: outdata = 32'd19097;
			46440: outdata = 32'd19096;
			46441: outdata = 32'd19095;
			46442: outdata = 32'd19094;
			46443: outdata = 32'd19093;
			46444: outdata = 32'd19092;
			46445: outdata = 32'd19091;
			46446: outdata = 32'd19090;
			46447: outdata = 32'd19089;
			46448: outdata = 32'd19088;
			46449: outdata = 32'd19087;
			46450: outdata = 32'd19086;
			46451: outdata = 32'd19085;
			46452: outdata = 32'd19084;
			46453: outdata = 32'd19083;
			46454: outdata = 32'd19082;
			46455: outdata = 32'd19081;
			46456: outdata = 32'd19080;
			46457: outdata = 32'd19079;
			46458: outdata = 32'd19078;
			46459: outdata = 32'd19077;
			46460: outdata = 32'd19076;
			46461: outdata = 32'd19075;
			46462: outdata = 32'd19074;
			46463: outdata = 32'd19073;
			46464: outdata = 32'd19072;
			46465: outdata = 32'd19071;
			46466: outdata = 32'd19070;
			46467: outdata = 32'd19069;
			46468: outdata = 32'd19068;
			46469: outdata = 32'd19067;
			46470: outdata = 32'd19066;
			46471: outdata = 32'd19065;
			46472: outdata = 32'd19064;
			46473: outdata = 32'd19063;
			46474: outdata = 32'd19062;
			46475: outdata = 32'd19061;
			46476: outdata = 32'd19060;
			46477: outdata = 32'd19059;
			46478: outdata = 32'd19058;
			46479: outdata = 32'd19057;
			46480: outdata = 32'd19056;
			46481: outdata = 32'd19055;
			46482: outdata = 32'd19054;
			46483: outdata = 32'd19053;
			46484: outdata = 32'd19052;
			46485: outdata = 32'd19051;
			46486: outdata = 32'd19050;
			46487: outdata = 32'd19049;
			46488: outdata = 32'd19048;
			46489: outdata = 32'd19047;
			46490: outdata = 32'd19046;
			46491: outdata = 32'd19045;
			46492: outdata = 32'd19044;
			46493: outdata = 32'd19043;
			46494: outdata = 32'd19042;
			46495: outdata = 32'd19041;
			46496: outdata = 32'd19040;
			46497: outdata = 32'd19039;
			46498: outdata = 32'd19038;
			46499: outdata = 32'd19037;
			46500: outdata = 32'd19036;
			46501: outdata = 32'd19035;
			46502: outdata = 32'd19034;
			46503: outdata = 32'd19033;
			46504: outdata = 32'd19032;
			46505: outdata = 32'd19031;
			46506: outdata = 32'd19030;
			46507: outdata = 32'd19029;
			46508: outdata = 32'd19028;
			46509: outdata = 32'd19027;
			46510: outdata = 32'd19026;
			46511: outdata = 32'd19025;
			46512: outdata = 32'd19024;
			46513: outdata = 32'd19023;
			46514: outdata = 32'd19022;
			46515: outdata = 32'd19021;
			46516: outdata = 32'd19020;
			46517: outdata = 32'd19019;
			46518: outdata = 32'd19018;
			46519: outdata = 32'd19017;
			46520: outdata = 32'd19016;
			46521: outdata = 32'd19015;
			46522: outdata = 32'd19014;
			46523: outdata = 32'd19013;
			46524: outdata = 32'd19012;
			46525: outdata = 32'd19011;
			46526: outdata = 32'd19010;
			46527: outdata = 32'd19009;
			46528: outdata = 32'd19008;
			46529: outdata = 32'd19007;
			46530: outdata = 32'd19006;
			46531: outdata = 32'd19005;
			46532: outdata = 32'd19004;
			46533: outdata = 32'd19003;
			46534: outdata = 32'd19002;
			46535: outdata = 32'd19001;
			46536: outdata = 32'd19000;
			46537: outdata = 32'd18999;
			46538: outdata = 32'd18998;
			46539: outdata = 32'd18997;
			46540: outdata = 32'd18996;
			46541: outdata = 32'd18995;
			46542: outdata = 32'd18994;
			46543: outdata = 32'd18993;
			46544: outdata = 32'd18992;
			46545: outdata = 32'd18991;
			46546: outdata = 32'd18990;
			46547: outdata = 32'd18989;
			46548: outdata = 32'd18988;
			46549: outdata = 32'd18987;
			46550: outdata = 32'd18986;
			46551: outdata = 32'd18985;
			46552: outdata = 32'd18984;
			46553: outdata = 32'd18983;
			46554: outdata = 32'd18982;
			46555: outdata = 32'd18981;
			46556: outdata = 32'd18980;
			46557: outdata = 32'd18979;
			46558: outdata = 32'd18978;
			46559: outdata = 32'd18977;
			46560: outdata = 32'd18976;
			46561: outdata = 32'd18975;
			46562: outdata = 32'd18974;
			46563: outdata = 32'd18973;
			46564: outdata = 32'd18972;
			46565: outdata = 32'd18971;
			46566: outdata = 32'd18970;
			46567: outdata = 32'd18969;
			46568: outdata = 32'd18968;
			46569: outdata = 32'd18967;
			46570: outdata = 32'd18966;
			46571: outdata = 32'd18965;
			46572: outdata = 32'd18964;
			46573: outdata = 32'd18963;
			46574: outdata = 32'd18962;
			46575: outdata = 32'd18961;
			46576: outdata = 32'd18960;
			46577: outdata = 32'd18959;
			46578: outdata = 32'd18958;
			46579: outdata = 32'd18957;
			46580: outdata = 32'd18956;
			46581: outdata = 32'd18955;
			46582: outdata = 32'd18954;
			46583: outdata = 32'd18953;
			46584: outdata = 32'd18952;
			46585: outdata = 32'd18951;
			46586: outdata = 32'd18950;
			46587: outdata = 32'd18949;
			46588: outdata = 32'd18948;
			46589: outdata = 32'd18947;
			46590: outdata = 32'd18946;
			46591: outdata = 32'd18945;
			46592: outdata = 32'd18944;
			46593: outdata = 32'd18943;
			46594: outdata = 32'd18942;
			46595: outdata = 32'd18941;
			46596: outdata = 32'd18940;
			46597: outdata = 32'd18939;
			46598: outdata = 32'd18938;
			46599: outdata = 32'd18937;
			46600: outdata = 32'd18936;
			46601: outdata = 32'd18935;
			46602: outdata = 32'd18934;
			46603: outdata = 32'd18933;
			46604: outdata = 32'd18932;
			46605: outdata = 32'd18931;
			46606: outdata = 32'd18930;
			46607: outdata = 32'd18929;
			46608: outdata = 32'd18928;
			46609: outdata = 32'd18927;
			46610: outdata = 32'd18926;
			46611: outdata = 32'd18925;
			46612: outdata = 32'd18924;
			46613: outdata = 32'd18923;
			46614: outdata = 32'd18922;
			46615: outdata = 32'd18921;
			46616: outdata = 32'd18920;
			46617: outdata = 32'd18919;
			46618: outdata = 32'd18918;
			46619: outdata = 32'd18917;
			46620: outdata = 32'd18916;
			46621: outdata = 32'd18915;
			46622: outdata = 32'd18914;
			46623: outdata = 32'd18913;
			46624: outdata = 32'd18912;
			46625: outdata = 32'd18911;
			46626: outdata = 32'd18910;
			46627: outdata = 32'd18909;
			46628: outdata = 32'd18908;
			46629: outdata = 32'd18907;
			46630: outdata = 32'd18906;
			46631: outdata = 32'd18905;
			46632: outdata = 32'd18904;
			46633: outdata = 32'd18903;
			46634: outdata = 32'd18902;
			46635: outdata = 32'd18901;
			46636: outdata = 32'd18900;
			46637: outdata = 32'd18899;
			46638: outdata = 32'd18898;
			46639: outdata = 32'd18897;
			46640: outdata = 32'd18896;
			46641: outdata = 32'd18895;
			46642: outdata = 32'd18894;
			46643: outdata = 32'd18893;
			46644: outdata = 32'd18892;
			46645: outdata = 32'd18891;
			46646: outdata = 32'd18890;
			46647: outdata = 32'd18889;
			46648: outdata = 32'd18888;
			46649: outdata = 32'd18887;
			46650: outdata = 32'd18886;
			46651: outdata = 32'd18885;
			46652: outdata = 32'd18884;
			46653: outdata = 32'd18883;
			46654: outdata = 32'd18882;
			46655: outdata = 32'd18881;
			46656: outdata = 32'd18880;
			46657: outdata = 32'd18879;
			46658: outdata = 32'd18878;
			46659: outdata = 32'd18877;
			46660: outdata = 32'd18876;
			46661: outdata = 32'd18875;
			46662: outdata = 32'd18874;
			46663: outdata = 32'd18873;
			46664: outdata = 32'd18872;
			46665: outdata = 32'd18871;
			46666: outdata = 32'd18870;
			46667: outdata = 32'd18869;
			46668: outdata = 32'd18868;
			46669: outdata = 32'd18867;
			46670: outdata = 32'd18866;
			46671: outdata = 32'd18865;
			46672: outdata = 32'd18864;
			46673: outdata = 32'd18863;
			46674: outdata = 32'd18862;
			46675: outdata = 32'd18861;
			46676: outdata = 32'd18860;
			46677: outdata = 32'd18859;
			46678: outdata = 32'd18858;
			46679: outdata = 32'd18857;
			46680: outdata = 32'd18856;
			46681: outdata = 32'd18855;
			46682: outdata = 32'd18854;
			46683: outdata = 32'd18853;
			46684: outdata = 32'd18852;
			46685: outdata = 32'd18851;
			46686: outdata = 32'd18850;
			46687: outdata = 32'd18849;
			46688: outdata = 32'd18848;
			46689: outdata = 32'd18847;
			46690: outdata = 32'd18846;
			46691: outdata = 32'd18845;
			46692: outdata = 32'd18844;
			46693: outdata = 32'd18843;
			46694: outdata = 32'd18842;
			46695: outdata = 32'd18841;
			46696: outdata = 32'd18840;
			46697: outdata = 32'd18839;
			46698: outdata = 32'd18838;
			46699: outdata = 32'd18837;
			46700: outdata = 32'd18836;
			46701: outdata = 32'd18835;
			46702: outdata = 32'd18834;
			46703: outdata = 32'd18833;
			46704: outdata = 32'd18832;
			46705: outdata = 32'd18831;
			46706: outdata = 32'd18830;
			46707: outdata = 32'd18829;
			46708: outdata = 32'd18828;
			46709: outdata = 32'd18827;
			46710: outdata = 32'd18826;
			46711: outdata = 32'd18825;
			46712: outdata = 32'd18824;
			46713: outdata = 32'd18823;
			46714: outdata = 32'd18822;
			46715: outdata = 32'd18821;
			46716: outdata = 32'd18820;
			46717: outdata = 32'd18819;
			46718: outdata = 32'd18818;
			46719: outdata = 32'd18817;
			46720: outdata = 32'd18816;
			46721: outdata = 32'd18815;
			46722: outdata = 32'd18814;
			46723: outdata = 32'd18813;
			46724: outdata = 32'd18812;
			46725: outdata = 32'd18811;
			46726: outdata = 32'd18810;
			46727: outdata = 32'd18809;
			46728: outdata = 32'd18808;
			46729: outdata = 32'd18807;
			46730: outdata = 32'd18806;
			46731: outdata = 32'd18805;
			46732: outdata = 32'd18804;
			46733: outdata = 32'd18803;
			46734: outdata = 32'd18802;
			46735: outdata = 32'd18801;
			46736: outdata = 32'd18800;
			46737: outdata = 32'd18799;
			46738: outdata = 32'd18798;
			46739: outdata = 32'd18797;
			46740: outdata = 32'd18796;
			46741: outdata = 32'd18795;
			46742: outdata = 32'd18794;
			46743: outdata = 32'd18793;
			46744: outdata = 32'd18792;
			46745: outdata = 32'd18791;
			46746: outdata = 32'd18790;
			46747: outdata = 32'd18789;
			46748: outdata = 32'd18788;
			46749: outdata = 32'd18787;
			46750: outdata = 32'd18786;
			46751: outdata = 32'd18785;
			46752: outdata = 32'd18784;
			46753: outdata = 32'd18783;
			46754: outdata = 32'd18782;
			46755: outdata = 32'd18781;
			46756: outdata = 32'd18780;
			46757: outdata = 32'd18779;
			46758: outdata = 32'd18778;
			46759: outdata = 32'd18777;
			46760: outdata = 32'd18776;
			46761: outdata = 32'd18775;
			46762: outdata = 32'd18774;
			46763: outdata = 32'd18773;
			46764: outdata = 32'd18772;
			46765: outdata = 32'd18771;
			46766: outdata = 32'd18770;
			46767: outdata = 32'd18769;
			46768: outdata = 32'd18768;
			46769: outdata = 32'd18767;
			46770: outdata = 32'd18766;
			46771: outdata = 32'd18765;
			46772: outdata = 32'd18764;
			46773: outdata = 32'd18763;
			46774: outdata = 32'd18762;
			46775: outdata = 32'd18761;
			46776: outdata = 32'd18760;
			46777: outdata = 32'd18759;
			46778: outdata = 32'd18758;
			46779: outdata = 32'd18757;
			46780: outdata = 32'd18756;
			46781: outdata = 32'd18755;
			46782: outdata = 32'd18754;
			46783: outdata = 32'd18753;
			46784: outdata = 32'd18752;
			46785: outdata = 32'd18751;
			46786: outdata = 32'd18750;
			46787: outdata = 32'd18749;
			46788: outdata = 32'd18748;
			46789: outdata = 32'd18747;
			46790: outdata = 32'd18746;
			46791: outdata = 32'd18745;
			46792: outdata = 32'd18744;
			46793: outdata = 32'd18743;
			46794: outdata = 32'd18742;
			46795: outdata = 32'd18741;
			46796: outdata = 32'd18740;
			46797: outdata = 32'd18739;
			46798: outdata = 32'd18738;
			46799: outdata = 32'd18737;
			46800: outdata = 32'd18736;
			46801: outdata = 32'd18735;
			46802: outdata = 32'd18734;
			46803: outdata = 32'd18733;
			46804: outdata = 32'd18732;
			46805: outdata = 32'd18731;
			46806: outdata = 32'd18730;
			46807: outdata = 32'd18729;
			46808: outdata = 32'd18728;
			46809: outdata = 32'd18727;
			46810: outdata = 32'd18726;
			46811: outdata = 32'd18725;
			46812: outdata = 32'd18724;
			46813: outdata = 32'd18723;
			46814: outdata = 32'd18722;
			46815: outdata = 32'd18721;
			46816: outdata = 32'd18720;
			46817: outdata = 32'd18719;
			46818: outdata = 32'd18718;
			46819: outdata = 32'd18717;
			46820: outdata = 32'd18716;
			46821: outdata = 32'd18715;
			46822: outdata = 32'd18714;
			46823: outdata = 32'd18713;
			46824: outdata = 32'd18712;
			46825: outdata = 32'd18711;
			46826: outdata = 32'd18710;
			46827: outdata = 32'd18709;
			46828: outdata = 32'd18708;
			46829: outdata = 32'd18707;
			46830: outdata = 32'd18706;
			46831: outdata = 32'd18705;
			46832: outdata = 32'd18704;
			46833: outdata = 32'd18703;
			46834: outdata = 32'd18702;
			46835: outdata = 32'd18701;
			46836: outdata = 32'd18700;
			46837: outdata = 32'd18699;
			46838: outdata = 32'd18698;
			46839: outdata = 32'd18697;
			46840: outdata = 32'd18696;
			46841: outdata = 32'd18695;
			46842: outdata = 32'd18694;
			46843: outdata = 32'd18693;
			46844: outdata = 32'd18692;
			46845: outdata = 32'd18691;
			46846: outdata = 32'd18690;
			46847: outdata = 32'd18689;
			46848: outdata = 32'd18688;
			46849: outdata = 32'd18687;
			46850: outdata = 32'd18686;
			46851: outdata = 32'd18685;
			46852: outdata = 32'd18684;
			46853: outdata = 32'd18683;
			46854: outdata = 32'd18682;
			46855: outdata = 32'd18681;
			46856: outdata = 32'd18680;
			46857: outdata = 32'd18679;
			46858: outdata = 32'd18678;
			46859: outdata = 32'd18677;
			46860: outdata = 32'd18676;
			46861: outdata = 32'd18675;
			46862: outdata = 32'd18674;
			46863: outdata = 32'd18673;
			46864: outdata = 32'd18672;
			46865: outdata = 32'd18671;
			46866: outdata = 32'd18670;
			46867: outdata = 32'd18669;
			46868: outdata = 32'd18668;
			46869: outdata = 32'd18667;
			46870: outdata = 32'd18666;
			46871: outdata = 32'd18665;
			46872: outdata = 32'd18664;
			46873: outdata = 32'd18663;
			46874: outdata = 32'd18662;
			46875: outdata = 32'd18661;
			46876: outdata = 32'd18660;
			46877: outdata = 32'd18659;
			46878: outdata = 32'd18658;
			46879: outdata = 32'd18657;
			46880: outdata = 32'd18656;
			46881: outdata = 32'd18655;
			46882: outdata = 32'd18654;
			46883: outdata = 32'd18653;
			46884: outdata = 32'd18652;
			46885: outdata = 32'd18651;
			46886: outdata = 32'd18650;
			46887: outdata = 32'd18649;
			46888: outdata = 32'd18648;
			46889: outdata = 32'd18647;
			46890: outdata = 32'd18646;
			46891: outdata = 32'd18645;
			46892: outdata = 32'd18644;
			46893: outdata = 32'd18643;
			46894: outdata = 32'd18642;
			46895: outdata = 32'd18641;
			46896: outdata = 32'd18640;
			46897: outdata = 32'd18639;
			46898: outdata = 32'd18638;
			46899: outdata = 32'd18637;
			46900: outdata = 32'd18636;
			46901: outdata = 32'd18635;
			46902: outdata = 32'd18634;
			46903: outdata = 32'd18633;
			46904: outdata = 32'd18632;
			46905: outdata = 32'd18631;
			46906: outdata = 32'd18630;
			46907: outdata = 32'd18629;
			46908: outdata = 32'd18628;
			46909: outdata = 32'd18627;
			46910: outdata = 32'd18626;
			46911: outdata = 32'd18625;
			46912: outdata = 32'd18624;
			46913: outdata = 32'd18623;
			46914: outdata = 32'd18622;
			46915: outdata = 32'd18621;
			46916: outdata = 32'd18620;
			46917: outdata = 32'd18619;
			46918: outdata = 32'd18618;
			46919: outdata = 32'd18617;
			46920: outdata = 32'd18616;
			46921: outdata = 32'd18615;
			46922: outdata = 32'd18614;
			46923: outdata = 32'd18613;
			46924: outdata = 32'd18612;
			46925: outdata = 32'd18611;
			46926: outdata = 32'd18610;
			46927: outdata = 32'd18609;
			46928: outdata = 32'd18608;
			46929: outdata = 32'd18607;
			46930: outdata = 32'd18606;
			46931: outdata = 32'd18605;
			46932: outdata = 32'd18604;
			46933: outdata = 32'd18603;
			46934: outdata = 32'd18602;
			46935: outdata = 32'd18601;
			46936: outdata = 32'd18600;
			46937: outdata = 32'd18599;
			46938: outdata = 32'd18598;
			46939: outdata = 32'd18597;
			46940: outdata = 32'd18596;
			46941: outdata = 32'd18595;
			46942: outdata = 32'd18594;
			46943: outdata = 32'd18593;
			46944: outdata = 32'd18592;
			46945: outdata = 32'd18591;
			46946: outdata = 32'd18590;
			46947: outdata = 32'd18589;
			46948: outdata = 32'd18588;
			46949: outdata = 32'd18587;
			46950: outdata = 32'd18586;
			46951: outdata = 32'd18585;
			46952: outdata = 32'd18584;
			46953: outdata = 32'd18583;
			46954: outdata = 32'd18582;
			46955: outdata = 32'd18581;
			46956: outdata = 32'd18580;
			46957: outdata = 32'd18579;
			46958: outdata = 32'd18578;
			46959: outdata = 32'd18577;
			46960: outdata = 32'd18576;
			46961: outdata = 32'd18575;
			46962: outdata = 32'd18574;
			46963: outdata = 32'd18573;
			46964: outdata = 32'd18572;
			46965: outdata = 32'd18571;
			46966: outdata = 32'd18570;
			46967: outdata = 32'd18569;
			46968: outdata = 32'd18568;
			46969: outdata = 32'd18567;
			46970: outdata = 32'd18566;
			46971: outdata = 32'd18565;
			46972: outdata = 32'd18564;
			46973: outdata = 32'd18563;
			46974: outdata = 32'd18562;
			46975: outdata = 32'd18561;
			46976: outdata = 32'd18560;
			46977: outdata = 32'd18559;
			46978: outdata = 32'd18558;
			46979: outdata = 32'd18557;
			46980: outdata = 32'd18556;
			46981: outdata = 32'd18555;
			46982: outdata = 32'd18554;
			46983: outdata = 32'd18553;
			46984: outdata = 32'd18552;
			46985: outdata = 32'd18551;
			46986: outdata = 32'd18550;
			46987: outdata = 32'd18549;
			46988: outdata = 32'd18548;
			46989: outdata = 32'd18547;
			46990: outdata = 32'd18546;
			46991: outdata = 32'd18545;
			46992: outdata = 32'd18544;
			46993: outdata = 32'd18543;
			46994: outdata = 32'd18542;
			46995: outdata = 32'd18541;
			46996: outdata = 32'd18540;
			46997: outdata = 32'd18539;
			46998: outdata = 32'd18538;
			46999: outdata = 32'd18537;
			47000: outdata = 32'd18536;
			47001: outdata = 32'd18535;
			47002: outdata = 32'd18534;
			47003: outdata = 32'd18533;
			47004: outdata = 32'd18532;
			47005: outdata = 32'd18531;
			47006: outdata = 32'd18530;
			47007: outdata = 32'd18529;
			47008: outdata = 32'd18528;
			47009: outdata = 32'd18527;
			47010: outdata = 32'd18526;
			47011: outdata = 32'd18525;
			47012: outdata = 32'd18524;
			47013: outdata = 32'd18523;
			47014: outdata = 32'd18522;
			47015: outdata = 32'd18521;
			47016: outdata = 32'd18520;
			47017: outdata = 32'd18519;
			47018: outdata = 32'd18518;
			47019: outdata = 32'd18517;
			47020: outdata = 32'd18516;
			47021: outdata = 32'd18515;
			47022: outdata = 32'd18514;
			47023: outdata = 32'd18513;
			47024: outdata = 32'd18512;
			47025: outdata = 32'd18511;
			47026: outdata = 32'd18510;
			47027: outdata = 32'd18509;
			47028: outdata = 32'd18508;
			47029: outdata = 32'd18507;
			47030: outdata = 32'd18506;
			47031: outdata = 32'd18505;
			47032: outdata = 32'd18504;
			47033: outdata = 32'd18503;
			47034: outdata = 32'd18502;
			47035: outdata = 32'd18501;
			47036: outdata = 32'd18500;
			47037: outdata = 32'd18499;
			47038: outdata = 32'd18498;
			47039: outdata = 32'd18497;
			47040: outdata = 32'd18496;
			47041: outdata = 32'd18495;
			47042: outdata = 32'd18494;
			47043: outdata = 32'd18493;
			47044: outdata = 32'd18492;
			47045: outdata = 32'd18491;
			47046: outdata = 32'd18490;
			47047: outdata = 32'd18489;
			47048: outdata = 32'd18488;
			47049: outdata = 32'd18487;
			47050: outdata = 32'd18486;
			47051: outdata = 32'd18485;
			47052: outdata = 32'd18484;
			47053: outdata = 32'd18483;
			47054: outdata = 32'd18482;
			47055: outdata = 32'd18481;
			47056: outdata = 32'd18480;
			47057: outdata = 32'd18479;
			47058: outdata = 32'd18478;
			47059: outdata = 32'd18477;
			47060: outdata = 32'd18476;
			47061: outdata = 32'd18475;
			47062: outdata = 32'd18474;
			47063: outdata = 32'd18473;
			47064: outdata = 32'd18472;
			47065: outdata = 32'd18471;
			47066: outdata = 32'd18470;
			47067: outdata = 32'd18469;
			47068: outdata = 32'd18468;
			47069: outdata = 32'd18467;
			47070: outdata = 32'd18466;
			47071: outdata = 32'd18465;
			47072: outdata = 32'd18464;
			47073: outdata = 32'd18463;
			47074: outdata = 32'd18462;
			47075: outdata = 32'd18461;
			47076: outdata = 32'd18460;
			47077: outdata = 32'd18459;
			47078: outdata = 32'd18458;
			47079: outdata = 32'd18457;
			47080: outdata = 32'd18456;
			47081: outdata = 32'd18455;
			47082: outdata = 32'd18454;
			47083: outdata = 32'd18453;
			47084: outdata = 32'd18452;
			47085: outdata = 32'd18451;
			47086: outdata = 32'd18450;
			47087: outdata = 32'd18449;
			47088: outdata = 32'd18448;
			47089: outdata = 32'd18447;
			47090: outdata = 32'd18446;
			47091: outdata = 32'd18445;
			47092: outdata = 32'd18444;
			47093: outdata = 32'd18443;
			47094: outdata = 32'd18442;
			47095: outdata = 32'd18441;
			47096: outdata = 32'd18440;
			47097: outdata = 32'd18439;
			47098: outdata = 32'd18438;
			47099: outdata = 32'd18437;
			47100: outdata = 32'd18436;
			47101: outdata = 32'd18435;
			47102: outdata = 32'd18434;
			47103: outdata = 32'd18433;
			47104: outdata = 32'd18432;
			47105: outdata = 32'd18431;
			47106: outdata = 32'd18430;
			47107: outdata = 32'd18429;
			47108: outdata = 32'd18428;
			47109: outdata = 32'd18427;
			47110: outdata = 32'd18426;
			47111: outdata = 32'd18425;
			47112: outdata = 32'd18424;
			47113: outdata = 32'd18423;
			47114: outdata = 32'd18422;
			47115: outdata = 32'd18421;
			47116: outdata = 32'd18420;
			47117: outdata = 32'd18419;
			47118: outdata = 32'd18418;
			47119: outdata = 32'd18417;
			47120: outdata = 32'd18416;
			47121: outdata = 32'd18415;
			47122: outdata = 32'd18414;
			47123: outdata = 32'd18413;
			47124: outdata = 32'd18412;
			47125: outdata = 32'd18411;
			47126: outdata = 32'd18410;
			47127: outdata = 32'd18409;
			47128: outdata = 32'd18408;
			47129: outdata = 32'd18407;
			47130: outdata = 32'd18406;
			47131: outdata = 32'd18405;
			47132: outdata = 32'd18404;
			47133: outdata = 32'd18403;
			47134: outdata = 32'd18402;
			47135: outdata = 32'd18401;
			47136: outdata = 32'd18400;
			47137: outdata = 32'd18399;
			47138: outdata = 32'd18398;
			47139: outdata = 32'd18397;
			47140: outdata = 32'd18396;
			47141: outdata = 32'd18395;
			47142: outdata = 32'd18394;
			47143: outdata = 32'd18393;
			47144: outdata = 32'd18392;
			47145: outdata = 32'd18391;
			47146: outdata = 32'd18390;
			47147: outdata = 32'd18389;
			47148: outdata = 32'd18388;
			47149: outdata = 32'd18387;
			47150: outdata = 32'd18386;
			47151: outdata = 32'd18385;
			47152: outdata = 32'd18384;
			47153: outdata = 32'd18383;
			47154: outdata = 32'd18382;
			47155: outdata = 32'd18381;
			47156: outdata = 32'd18380;
			47157: outdata = 32'd18379;
			47158: outdata = 32'd18378;
			47159: outdata = 32'd18377;
			47160: outdata = 32'd18376;
			47161: outdata = 32'd18375;
			47162: outdata = 32'd18374;
			47163: outdata = 32'd18373;
			47164: outdata = 32'd18372;
			47165: outdata = 32'd18371;
			47166: outdata = 32'd18370;
			47167: outdata = 32'd18369;
			47168: outdata = 32'd18368;
			47169: outdata = 32'd18367;
			47170: outdata = 32'd18366;
			47171: outdata = 32'd18365;
			47172: outdata = 32'd18364;
			47173: outdata = 32'd18363;
			47174: outdata = 32'd18362;
			47175: outdata = 32'd18361;
			47176: outdata = 32'd18360;
			47177: outdata = 32'd18359;
			47178: outdata = 32'd18358;
			47179: outdata = 32'd18357;
			47180: outdata = 32'd18356;
			47181: outdata = 32'd18355;
			47182: outdata = 32'd18354;
			47183: outdata = 32'd18353;
			47184: outdata = 32'd18352;
			47185: outdata = 32'd18351;
			47186: outdata = 32'd18350;
			47187: outdata = 32'd18349;
			47188: outdata = 32'd18348;
			47189: outdata = 32'd18347;
			47190: outdata = 32'd18346;
			47191: outdata = 32'd18345;
			47192: outdata = 32'd18344;
			47193: outdata = 32'd18343;
			47194: outdata = 32'd18342;
			47195: outdata = 32'd18341;
			47196: outdata = 32'd18340;
			47197: outdata = 32'd18339;
			47198: outdata = 32'd18338;
			47199: outdata = 32'd18337;
			47200: outdata = 32'd18336;
			47201: outdata = 32'd18335;
			47202: outdata = 32'd18334;
			47203: outdata = 32'd18333;
			47204: outdata = 32'd18332;
			47205: outdata = 32'd18331;
			47206: outdata = 32'd18330;
			47207: outdata = 32'd18329;
			47208: outdata = 32'd18328;
			47209: outdata = 32'd18327;
			47210: outdata = 32'd18326;
			47211: outdata = 32'd18325;
			47212: outdata = 32'd18324;
			47213: outdata = 32'd18323;
			47214: outdata = 32'd18322;
			47215: outdata = 32'd18321;
			47216: outdata = 32'd18320;
			47217: outdata = 32'd18319;
			47218: outdata = 32'd18318;
			47219: outdata = 32'd18317;
			47220: outdata = 32'd18316;
			47221: outdata = 32'd18315;
			47222: outdata = 32'd18314;
			47223: outdata = 32'd18313;
			47224: outdata = 32'd18312;
			47225: outdata = 32'd18311;
			47226: outdata = 32'd18310;
			47227: outdata = 32'd18309;
			47228: outdata = 32'd18308;
			47229: outdata = 32'd18307;
			47230: outdata = 32'd18306;
			47231: outdata = 32'd18305;
			47232: outdata = 32'd18304;
			47233: outdata = 32'd18303;
			47234: outdata = 32'd18302;
			47235: outdata = 32'd18301;
			47236: outdata = 32'd18300;
			47237: outdata = 32'd18299;
			47238: outdata = 32'd18298;
			47239: outdata = 32'd18297;
			47240: outdata = 32'd18296;
			47241: outdata = 32'd18295;
			47242: outdata = 32'd18294;
			47243: outdata = 32'd18293;
			47244: outdata = 32'd18292;
			47245: outdata = 32'd18291;
			47246: outdata = 32'd18290;
			47247: outdata = 32'd18289;
			47248: outdata = 32'd18288;
			47249: outdata = 32'd18287;
			47250: outdata = 32'd18286;
			47251: outdata = 32'd18285;
			47252: outdata = 32'd18284;
			47253: outdata = 32'd18283;
			47254: outdata = 32'd18282;
			47255: outdata = 32'd18281;
			47256: outdata = 32'd18280;
			47257: outdata = 32'd18279;
			47258: outdata = 32'd18278;
			47259: outdata = 32'd18277;
			47260: outdata = 32'd18276;
			47261: outdata = 32'd18275;
			47262: outdata = 32'd18274;
			47263: outdata = 32'd18273;
			47264: outdata = 32'd18272;
			47265: outdata = 32'd18271;
			47266: outdata = 32'd18270;
			47267: outdata = 32'd18269;
			47268: outdata = 32'd18268;
			47269: outdata = 32'd18267;
			47270: outdata = 32'd18266;
			47271: outdata = 32'd18265;
			47272: outdata = 32'd18264;
			47273: outdata = 32'd18263;
			47274: outdata = 32'd18262;
			47275: outdata = 32'd18261;
			47276: outdata = 32'd18260;
			47277: outdata = 32'd18259;
			47278: outdata = 32'd18258;
			47279: outdata = 32'd18257;
			47280: outdata = 32'd18256;
			47281: outdata = 32'd18255;
			47282: outdata = 32'd18254;
			47283: outdata = 32'd18253;
			47284: outdata = 32'd18252;
			47285: outdata = 32'd18251;
			47286: outdata = 32'd18250;
			47287: outdata = 32'd18249;
			47288: outdata = 32'd18248;
			47289: outdata = 32'd18247;
			47290: outdata = 32'd18246;
			47291: outdata = 32'd18245;
			47292: outdata = 32'd18244;
			47293: outdata = 32'd18243;
			47294: outdata = 32'd18242;
			47295: outdata = 32'd18241;
			47296: outdata = 32'd18240;
			47297: outdata = 32'd18239;
			47298: outdata = 32'd18238;
			47299: outdata = 32'd18237;
			47300: outdata = 32'd18236;
			47301: outdata = 32'd18235;
			47302: outdata = 32'd18234;
			47303: outdata = 32'd18233;
			47304: outdata = 32'd18232;
			47305: outdata = 32'd18231;
			47306: outdata = 32'd18230;
			47307: outdata = 32'd18229;
			47308: outdata = 32'd18228;
			47309: outdata = 32'd18227;
			47310: outdata = 32'd18226;
			47311: outdata = 32'd18225;
			47312: outdata = 32'd18224;
			47313: outdata = 32'd18223;
			47314: outdata = 32'd18222;
			47315: outdata = 32'd18221;
			47316: outdata = 32'd18220;
			47317: outdata = 32'd18219;
			47318: outdata = 32'd18218;
			47319: outdata = 32'd18217;
			47320: outdata = 32'd18216;
			47321: outdata = 32'd18215;
			47322: outdata = 32'd18214;
			47323: outdata = 32'd18213;
			47324: outdata = 32'd18212;
			47325: outdata = 32'd18211;
			47326: outdata = 32'd18210;
			47327: outdata = 32'd18209;
			47328: outdata = 32'd18208;
			47329: outdata = 32'd18207;
			47330: outdata = 32'd18206;
			47331: outdata = 32'd18205;
			47332: outdata = 32'd18204;
			47333: outdata = 32'd18203;
			47334: outdata = 32'd18202;
			47335: outdata = 32'd18201;
			47336: outdata = 32'd18200;
			47337: outdata = 32'd18199;
			47338: outdata = 32'd18198;
			47339: outdata = 32'd18197;
			47340: outdata = 32'd18196;
			47341: outdata = 32'd18195;
			47342: outdata = 32'd18194;
			47343: outdata = 32'd18193;
			47344: outdata = 32'd18192;
			47345: outdata = 32'd18191;
			47346: outdata = 32'd18190;
			47347: outdata = 32'd18189;
			47348: outdata = 32'd18188;
			47349: outdata = 32'd18187;
			47350: outdata = 32'd18186;
			47351: outdata = 32'd18185;
			47352: outdata = 32'd18184;
			47353: outdata = 32'd18183;
			47354: outdata = 32'd18182;
			47355: outdata = 32'd18181;
			47356: outdata = 32'd18180;
			47357: outdata = 32'd18179;
			47358: outdata = 32'd18178;
			47359: outdata = 32'd18177;
			47360: outdata = 32'd18176;
			47361: outdata = 32'd18175;
			47362: outdata = 32'd18174;
			47363: outdata = 32'd18173;
			47364: outdata = 32'd18172;
			47365: outdata = 32'd18171;
			47366: outdata = 32'd18170;
			47367: outdata = 32'd18169;
			47368: outdata = 32'd18168;
			47369: outdata = 32'd18167;
			47370: outdata = 32'd18166;
			47371: outdata = 32'd18165;
			47372: outdata = 32'd18164;
			47373: outdata = 32'd18163;
			47374: outdata = 32'd18162;
			47375: outdata = 32'd18161;
			47376: outdata = 32'd18160;
			47377: outdata = 32'd18159;
			47378: outdata = 32'd18158;
			47379: outdata = 32'd18157;
			47380: outdata = 32'd18156;
			47381: outdata = 32'd18155;
			47382: outdata = 32'd18154;
			47383: outdata = 32'd18153;
			47384: outdata = 32'd18152;
			47385: outdata = 32'd18151;
			47386: outdata = 32'd18150;
			47387: outdata = 32'd18149;
			47388: outdata = 32'd18148;
			47389: outdata = 32'd18147;
			47390: outdata = 32'd18146;
			47391: outdata = 32'd18145;
			47392: outdata = 32'd18144;
			47393: outdata = 32'd18143;
			47394: outdata = 32'd18142;
			47395: outdata = 32'd18141;
			47396: outdata = 32'd18140;
			47397: outdata = 32'd18139;
			47398: outdata = 32'd18138;
			47399: outdata = 32'd18137;
			47400: outdata = 32'd18136;
			47401: outdata = 32'd18135;
			47402: outdata = 32'd18134;
			47403: outdata = 32'd18133;
			47404: outdata = 32'd18132;
			47405: outdata = 32'd18131;
			47406: outdata = 32'd18130;
			47407: outdata = 32'd18129;
			47408: outdata = 32'd18128;
			47409: outdata = 32'd18127;
			47410: outdata = 32'd18126;
			47411: outdata = 32'd18125;
			47412: outdata = 32'd18124;
			47413: outdata = 32'd18123;
			47414: outdata = 32'd18122;
			47415: outdata = 32'd18121;
			47416: outdata = 32'd18120;
			47417: outdata = 32'd18119;
			47418: outdata = 32'd18118;
			47419: outdata = 32'd18117;
			47420: outdata = 32'd18116;
			47421: outdata = 32'd18115;
			47422: outdata = 32'd18114;
			47423: outdata = 32'd18113;
			47424: outdata = 32'd18112;
			47425: outdata = 32'd18111;
			47426: outdata = 32'd18110;
			47427: outdata = 32'd18109;
			47428: outdata = 32'd18108;
			47429: outdata = 32'd18107;
			47430: outdata = 32'd18106;
			47431: outdata = 32'd18105;
			47432: outdata = 32'd18104;
			47433: outdata = 32'd18103;
			47434: outdata = 32'd18102;
			47435: outdata = 32'd18101;
			47436: outdata = 32'd18100;
			47437: outdata = 32'd18099;
			47438: outdata = 32'd18098;
			47439: outdata = 32'd18097;
			47440: outdata = 32'd18096;
			47441: outdata = 32'd18095;
			47442: outdata = 32'd18094;
			47443: outdata = 32'd18093;
			47444: outdata = 32'd18092;
			47445: outdata = 32'd18091;
			47446: outdata = 32'd18090;
			47447: outdata = 32'd18089;
			47448: outdata = 32'd18088;
			47449: outdata = 32'd18087;
			47450: outdata = 32'd18086;
			47451: outdata = 32'd18085;
			47452: outdata = 32'd18084;
			47453: outdata = 32'd18083;
			47454: outdata = 32'd18082;
			47455: outdata = 32'd18081;
			47456: outdata = 32'd18080;
			47457: outdata = 32'd18079;
			47458: outdata = 32'd18078;
			47459: outdata = 32'd18077;
			47460: outdata = 32'd18076;
			47461: outdata = 32'd18075;
			47462: outdata = 32'd18074;
			47463: outdata = 32'd18073;
			47464: outdata = 32'd18072;
			47465: outdata = 32'd18071;
			47466: outdata = 32'd18070;
			47467: outdata = 32'd18069;
			47468: outdata = 32'd18068;
			47469: outdata = 32'd18067;
			47470: outdata = 32'd18066;
			47471: outdata = 32'd18065;
			47472: outdata = 32'd18064;
			47473: outdata = 32'd18063;
			47474: outdata = 32'd18062;
			47475: outdata = 32'd18061;
			47476: outdata = 32'd18060;
			47477: outdata = 32'd18059;
			47478: outdata = 32'd18058;
			47479: outdata = 32'd18057;
			47480: outdata = 32'd18056;
			47481: outdata = 32'd18055;
			47482: outdata = 32'd18054;
			47483: outdata = 32'd18053;
			47484: outdata = 32'd18052;
			47485: outdata = 32'd18051;
			47486: outdata = 32'd18050;
			47487: outdata = 32'd18049;
			47488: outdata = 32'd18048;
			47489: outdata = 32'd18047;
			47490: outdata = 32'd18046;
			47491: outdata = 32'd18045;
			47492: outdata = 32'd18044;
			47493: outdata = 32'd18043;
			47494: outdata = 32'd18042;
			47495: outdata = 32'd18041;
			47496: outdata = 32'd18040;
			47497: outdata = 32'd18039;
			47498: outdata = 32'd18038;
			47499: outdata = 32'd18037;
			47500: outdata = 32'd18036;
			47501: outdata = 32'd18035;
			47502: outdata = 32'd18034;
			47503: outdata = 32'd18033;
			47504: outdata = 32'd18032;
			47505: outdata = 32'd18031;
			47506: outdata = 32'd18030;
			47507: outdata = 32'd18029;
			47508: outdata = 32'd18028;
			47509: outdata = 32'd18027;
			47510: outdata = 32'd18026;
			47511: outdata = 32'd18025;
			47512: outdata = 32'd18024;
			47513: outdata = 32'd18023;
			47514: outdata = 32'd18022;
			47515: outdata = 32'd18021;
			47516: outdata = 32'd18020;
			47517: outdata = 32'd18019;
			47518: outdata = 32'd18018;
			47519: outdata = 32'd18017;
			47520: outdata = 32'd18016;
			47521: outdata = 32'd18015;
			47522: outdata = 32'd18014;
			47523: outdata = 32'd18013;
			47524: outdata = 32'd18012;
			47525: outdata = 32'd18011;
			47526: outdata = 32'd18010;
			47527: outdata = 32'd18009;
			47528: outdata = 32'd18008;
			47529: outdata = 32'd18007;
			47530: outdata = 32'd18006;
			47531: outdata = 32'd18005;
			47532: outdata = 32'd18004;
			47533: outdata = 32'd18003;
			47534: outdata = 32'd18002;
			47535: outdata = 32'd18001;
			47536: outdata = 32'd18000;
			47537: outdata = 32'd17999;
			47538: outdata = 32'd17998;
			47539: outdata = 32'd17997;
			47540: outdata = 32'd17996;
			47541: outdata = 32'd17995;
			47542: outdata = 32'd17994;
			47543: outdata = 32'd17993;
			47544: outdata = 32'd17992;
			47545: outdata = 32'd17991;
			47546: outdata = 32'd17990;
			47547: outdata = 32'd17989;
			47548: outdata = 32'd17988;
			47549: outdata = 32'd17987;
			47550: outdata = 32'd17986;
			47551: outdata = 32'd17985;
			47552: outdata = 32'd17984;
			47553: outdata = 32'd17983;
			47554: outdata = 32'd17982;
			47555: outdata = 32'd17981;
			47556: outdata = 32'd17980;
			47557: outdata = 32'd17979;
			47558: outdata = 32'd17978;
			47559: outdata = 32'd17977;
			47560: outdata = 32'd17976;
			47561: outdata = 32'd17975;
			47562: outdata = 32'd17974;
			47563: outdata = 32'd17973;
			47564: outdata = 32'd17972;
			47565: outdata = 32'd17971;
			47566: outdata = 32'd17970;
			47567: outdata = 32'd17969;
			47568: outdata = 32'd17968;
			47569: outdata = 32'd17967;
			47570: outdata = 32'd17966;
			47571: outdata = 32'd17965;
			47572: outdata = 32'd17964;
			47573: outdata = 32'd17963;
			47574: outdata = 32'd17962;
			47575: outdata = 32'd17961;
			47576: outdata = 32'd17960;
			47577: outdata = 32'd17959;
			47578: outdata = 32'd17958;
			47579: outdata = 32'd17957;
			47580: outdata = 32'd17956;
			47581: outdata = 32'd17955;
			47582: outdata = 32'd17954;
			47583: outdata = 32'd17953;
			47584: outdata = 32'd17952;
			47585: outdata = 32'd17951;
			47586: outdata = 32'd17950;
			47587: outdata = 32'd17949;
			47588: outdata = 32'd17948;
			47589: outdata = 32'd17947;
			47590: outdata = 32'd17946;
			47591: outdata = 32'd17945;
			47592: outdata = 32'd17944;
			47593: outdata = 32'd17943;
			47594: outdata = 32'd17942;
			47595: outdata = 32'd17941;
			47596: outdata = 32'd17940;
			47597: outdata = 32'd17939;
			47598: outdata = 32'd17938;
			47599: outdata = 32'd17937;
			47600: outdata = 32'd17936;
			47601: outdata = 32'd17935;
			47602: outdata = 32'd17934;
			47603: outdata = 32'd17933;
			47604: outdata = 32'd17932;
			47605: outdata = 32'd17931;
			47606: outdata = 32'd17930;
			47607: outdata = 32'd17929;
			47608: outdata = 32'd17928;
			47609: outdata = 32'd17927;
			47610: outdata = 32'd17926;
			47611: outdata = 32'd17925;
			47612: outdata = 32'd17924;
			47613: outdata = 32'd17923;
			47614: outdata = 32'd17922;
			47615: outdata = 32'd17921;
			47616: outdata = 32'd17920;
			47617: outdata = 32'd17919;
			47618: outdata = 32'd17918;
			47619: outdata = 32'd17917;
			47620: outdata = 32'd17916;
			47621: outdata = 32'd17915;
			47622: outdata = 32'd17914;
			47623: outdata = 32'd17913;
			47624: outdata = 32'd17912;
			47625: outdata = 32'd17911;
			47626: outdata = 32'd17910;
			47627: outdata = 32'd17909;
			47628: outdata = 32'd17908;
			47629: outdata = 32'd17907;
			47630: outdata = 32'd17906;
			47631: outdata = 32'd17905;
			47632: outdata = 32'd17904;
			47633: outdata = 32'd17903;
			47634: outdata = 32'd17902;
			47635: outdata = 32'd17901;
			47636: outdata = 32'd17900;
			47637: outdata = 32'd17899;
			47638: outdata = 32'd17898;
			47639: outdata = 32'd17897;
			47640: outdata = 32'd17896;
			47641: outdata = 32'd17895;
			47642: outdata = 32'd17894;
			47643: outdata = 32'd17893;
			47644: outdata = 32'd17892;
			47645: outdata = 32'd17891;
			47646: outdata = 32'd17890;
			47647: outdata = 32'd17889;
			47648: outdata = 32'd17888;
			47649: outdata = 32'd17887;
			47650: outdata = 32'd17886;
			47651: outdata = 32'd17885;
			47652: outdata = 32'd17884;
			47653: outdata = 32'd17883;
			47654: outdata = 32'd17882;
			47655: outdata = 32'd17881;
			47656: outdata = 32'd17880;
			47657: outdata = 32'd17879;
			47658: outdata = 32'd17878;
			47659: outdata = 32'd17877;
			47660: outdata = 32'd17876;
			47661: outdata = 32'd17875;
			47662: outdata = 32'd17874;
			47663: outdata = 32'd17873;
			47664: outdata = 32'd17872;
			47665: outdata = 32'd17871;
			47666: outdata = 32'd17870;
			47667: outdata = 32'd17869;
			47668: outdata = 32'd17868;
			47669: outdata = 32'd17867;
			47670: outdata = 32'd17866;
			47671: outdata = 32'd17865;
			47672: outdata = 32'd17864;
			47673: outdata = 32'd17863;
			47674: outdata = 32'd17862;
			47675: outdata = 32'd17861;
			47676: outdata = 32'd17860;
			47677: outdata = 32'd17859;
			47678: outdata = 32'd17858;
			47679: outdata = 32'd17857;
			47680: outdata = 32'd17856;
			47681: outdata = 32'd17855;
			47682: outdata = 32'd17854;
			47683: outdata = 32'd17853;
			47684: outdata = 32'd17852;
			47685: outdata = 32'd17851;
			47686: outdata = 32'd17850;
			47687: outdata = 32'd17849;
			47688: outdata = 32'd17848;
			47689: outdata = 32'd17847;
			47690: outdata = 32'd17846;
			47691: outdata = 32'd17845;
			47692: outdata = 32'd17844;
			47693: outdata = 32'd17843;
			47694: outdata = 32'd17842;
			47695: outdata = 32'd17841;
			47696: outdata = 32'd17840;
			47697: outdata = 32'd17839;
			47698: outdata = 32'd17838;
			47699: outdata = 32'd17837;
			47700: outdata = 32'd17836;
			47701: outdata = 32'd17835;
			47702: outdata = 32'd17834;
			47703: outdata = 32'd17833;
			47704: outdata = 32'd17832;
			47705: outdata = 32'd17831;
			47706: outdata = 32'd17830;
			47707: outdata = 32'd17829;
			47708: outdata = 32'd17828;
			47709: outdata = 32'd17827;
			47710: outdata = 32'd17826;
			47711: outdata = 32'd17825;
			47712: outdata = 32'd17824;
			47713: outdata = 32'd17823;
			47714: outdata = 32'd17822;
			47715: outdata = 32'd17821;
			47716: outdata = 32'd17820;
			47717: outdata = 32'd17819;
			47718: outdata = 32'd17818;
			47719: outdata = 32'd17817;
			47720: outdata = 32'd17816;
			47721: outdata = 32'd17815;
			47722: outdata = 32'd17814;
			47723: outdata = 32'd17813;
			47724: outdata = 32'd17812;
			47725: outdata = 32'd17811;
			47726: outdata = 32'd17810;
			47727: outdata = 32'd17809;
			47728: outdata = 32'd17808;
			47729: outdata = 32'd17807;
			47730: outdata = 32'd17806;
			47731: outdata = 32'd17805;
			47732: outdata = 32'd17804;
			47733: outdata = 32'd17803;
			47734: outdata = 32'd17802;
			47735: outdata = 32'd17801;
			47736: outdata = 32'd17800;
			47737: outdata = 32'd17799;
			47738: outdata = 32'd17798;
			47739: outdata = 32'd17797;
			47740: outdata = 32'd17796;
			47741: outdata = 32'd17795;
			47742: outdata = 32'd17794;
			47743: outdata = 32'd17793;
			47744: outdata = 32'd17792;
			47745: outdata = 32'd17791;
			47746: outdata = 32'd17790;
			47747: outdata = 32'd17789;
			47748: outdata = 32'd17788;
			47749: outdata = 32'd17787;
			47750: outdata = 32'd17786;
			47751: outdata = 32'd17785;
			47752: outdata = 32'd17784;
			47753: outdata = 32'd17783;
			47754: outdata = 32'd17782;
			47755: outdata = 32'd17781;
			47756: outdata = 32'd17780;
			47757: outdata = 32'd17779;
			47758: outdata = 32'd17778;
			47759: outdata = 32'd17777;
			47760: outdata = 32'd17776;
			47761: outdata = 32'd17775;
			47762: outdata = 32'd17774;
			47763: outdata = 32'd17773;
			47764: outdata = 32'd17772;
			47765: outdata = 32'd17771;
			47766: outdata = 32'd17770;
			47767: outdata = 32'd17769;
			47768: outdata = 32'd17768;
			47769: outdata = 32'd17767;
			47770: outdata = 32'd17766;
			47771: outdata = 32'd17765;
			47772: outdata = 32'd17764;
			47773: outdata = 32'd17763;
			47774: outdata = 32'd17762;
			47775: outdata = 32'd17761;
			47776: outdata = 32'd17760;
			47777: outdata = 32'd17759;
			47778: outdata = 32'd17758;
			47779: outdata = 32'd17757;
			47780: outdata = 32'd17756;
			47781: outdata = 32'd17755;
			47782: outdata = 32'd17754;
			47783: outdata = 32'd17753;
			47784: outdata = 32'd17752;
			47785: outdata = 32'd17751;
			47786: outdata = 32'd17750;
			47787: outdata = 32'd17749;
			47788: outdata = 32'd17748;
			47789: outdata = 32'd17747;
			47790: outdata = 32'd17746;
			47791: outdata = 32'd17745;
			47792: outdata = 32'd17744;
			47793: outdata = 32'd17743;
			47794: outdata = 32'd17742;
			47795: outdata = 32'd17741;
			47796: outdata = 32'd17740;
			47797: outdata = 32'd17739;
			47798: outdata = 32'd17738;
			47799: outdata = 32'd17737;
			47800: outdata = 32'd17736;
			47801: outdata = 32'd17735;
			47802: outdata = 32'd17734;
			47803: outdata = 32'd17733;
			47804: outdata = 32'd17732;
			47805: outdata = 32'd17731;
			47806: outdata = 32'd17730;
			47807: outdata = 32'd17729;
			47808: outdata = 32'd17728;
			47809: outdata = 32'd17727;
			47810: outdata = 32'd17726;
			47811: outdata = 32'd17725;
			47812: outdata = 32'd17724;
			47813: outdata = 32'd17723;
			47814: outdata = 32'd17722;
			47815: outdata = 32'd17721;
			47816: outdata = 32'd17720;
			47817: outdata = 32'd17719;
			47818: outdata = 32'd17718;
			47819: outdata = 32'd17717;
			47820: outdata = 32'd17716;
			47821: outdata = 32'd17715;
			47822: outdata = 32'd17714;
			47823: outdata = 32'd17713;
			47824: outdata = 32'd17712;
			47825: outdata = 32'd17711;
			47826: outdata = 32'd17710;
			47827: outdata = 32'd17709;
			47828: outdata = 32'd17708;
			47829: outdata = 32'd17707;
			47830: outdata = 32'd17706;
			47831: outdata = 32'd17705;
			47832: outdata = 32'd17704;
			47833: outdata = 32'd17703;
			47834: outdata = 32'd17702;
			47835: outdata = 32'd17701;
			47836: outdata = 32'd17700;
			47837: outdata = 32'd17699;
			47838: outdata = 32'd17698;
			47839: outdata = 32'd17697;
			47840: outdata = 32'd17696;
			47841: outdata = 32'd17695;
			47842: outdata = 32'd17694;
			47843: outdata = 32'd17693;
			47844: outdata = 32'd17692;
			47845: outdata = 32'd17691;
			47846: outdata = 32'd17690;
			47847: outdata = 32'd17689;
			47848: outdata = 32'd17688;
			47849: outdata = 32'd17687;
			47850: outdata = 32'd17686;
			47851: outdata = 32'd17685;
			47852: outdata = 32'd17684;
			47853: outdata = 32'd17683;
			47854: outdata = 32'd17682;
			47855: outdata = 32'd17681;
			47856: outdata = 32'd17680;
			47857: outdata = 32'd17679;
			47858: outdata = 32'd17678;
			47859: outdata = 32'd17677;
			47860: outdata = 32'd17676;
			47861: outdata = 32'd17675;
			47862: outdata = 32'd17674;
			47863: outdata = 32'd17673;
			47864: outdata = 32'd17672;
			47865: outdata = 32'd17671;
			47866: outdata = 32'd17670;
			47867: outdata = 32'd17669;
			47868: outdata = 32'd17668;
			47869: outdata = 32'd17667;
			47870: outdata = 32'd17666;
			47871: outdata = 32'd17665;
			47872: outdata = 32'd17664;
			47873: outdata = 32'd17663;
			47874: outdata = 32'd17662;
			47875: outdata = 32'd17661;
			47876: outdata = 32'd17660;
			47877: outdata = 32'd17659;
			47878: outdata = 32'd17658;
			47879: outdata = 32'd17657;
			47880: outdata = 32'd17656;
			47881: outdata = 32'd17655;
			47882: outdata = 32'd17654;
			47883: outdata = 32'd17653;
			47884: outdata = 32'd17652;
			47885: outdata = 32'd17651;
			47886: outdata = 32'd17650;
			47887: outdata = 32'd17649;
			47888: outdata = 32'd17648;
			47889: outdata = 32'd17647;
			47890: outdata = 32'd17646;
			47891: outdata = 32'd17645;
			47892: outdata = 32'd17644;
			47893: outdata = 32'd17643;
			47894: outdata = 32'd17642;
			47895: outdata = 32'd17641;
			47896: outdata = 32'd17640;
			47897: outdata = 32'd17639;
			47898: outdata = 32'd17638;
			47899: outdata = 32'd17637;
			47900: outdata = 32'd17636;
			47901: outdata = 32'd17635;
			47902: outdata = 32'd17634;
			47903: outdata = 32'd17633;
			47904: outdata = 32'd17632;
			47905: outdata = 32'd17631;
			47906: outdata = 32'd17630;
			47907: outdata = 32'd17629;
			47908: outdata = 32'd17628;
			47909: outdata = 32'd17627;
			47910: outdata = 32'd17626;
			47911: outdata = 32'd17625;
			47912: outdata = 32'd17624;
			47913: outdata = 32'd17623;
			47914: outdata = 32'd17622;
			47915: outdata = 32'd17621;
			47916: outdata = 32'd17620;
			47917: outdata = 32'd17619;
			47918: outdata = 32'd17618;
			47919: outdata = 32'd17617;
			47920: outdata = 32'd17616;
			47921: outdata = 32'd17615;
			47922: outdata = 32'd17614;
			47923: outdata = 32'd17613;
			47924: outdata = 32'd17612;
			47925: outdata = 32'd17611;
			47926: outdata = 32'd17610;
			47927: outdata = 32'd17609;
			47928: outdata = 32'd17608;
			47929: outdata = 32'd17607;
			47930: outdata = 32'd17606;
			47931: outdata = 32'd17605;
			47932: outdata = 32'd17604;
			47933: outdata = 32'd17603;
			47934: outdata = 32'd17602;
			47935: outdata = 32'd17601;
			47936: outdata = 32'd17600;
			47937: outdata = 32'd17599;
			47938: outdata = 32'd17598;
			47939: outdata = 32'd17597;
			47940: outdata = 32'd17596;
			47941: outdata = 32'd17595;
			47942: outdata = 32'd17594;
			47943: outdata = 32'd17593;
			47944: outdata = 32'd17592;
			47945: outdata = 32'd17591;
			47946: outdata = 32'd17590;
			47947: outdata = 32'd17589;
			47948: outdata = 32'd17588;
			47949: outdata = 32'd17587;
			47950: outdata = 32'd17586;
			47951: outdata = 32'd17585;
			47952: outdata = 32'd17584;
			47953: outdata = 32'd17583;
			47954: outdata = 32'd17582;
			47955: outdata = 32'd17581;
			47956: outdata = 32'd17580;
			47957: outdata = 32'd17579;
			47958: outdata = 32'd17578;
			47959: outdata = 32'd17577;
			47960: outdata = 32'd17576;
			47961: outdata = 32'd17575;
			47962: outdata = 32'd17574;
			47963: outdata = 32'd17573;
			47964: outdata = 32'd17572;
			47965: outdata = 32'd17571;
			47966: outdata = 32'd17570;
			47967: outdata = 32'd17569;
			47968: outdata = 32'd17568;
			47969: outdata = 32'd17567;
			47970: outdata = 32'd17566;
			47971: outdata = 32'd17565;
			47972: outdata = 32'd17564;
			47973: outdata = 32'd17563;
			47974: outdata = 32'd17562;
			47975: outdata = 32'd17561;
			47976: outdata = 32'd17560;
			47977: outdata = 32'd17559;
			47978: outdata = 32'd17558;
			47979: outdata = 32'd17557;
			47980: outdata = 32'd17556;
			47981: outdata = 32'd17555;
			47982: outdata = 32'd17554;
			47983: outdata = 32'd17553;
			47984: outdata = 32'd17552;
			47985: outdata = 32'd17551;
			47986: outdata = 32'd17550;
			47987: outdata = 32'd17549;
			47988: outdata = 32'd17548;
			47989: outdata = 32'd17547;
			47990: outdata = 32'd17546;
			47991: outdata = 32'd17545;
			47992: outdata = 32'd17544;
			47993: outdata = 32'd17543;
			47994: outdata = 32'd17542;
			47995: outdata = 32'd17541;
			47996: outdata = 32'd17540;
			47997: outdata = 32'd17539;
			47998: outdata = 32'd17538;
			47999: outdata = 32'd17537;
			48000: outdata = 32'd17536;
			48001: outdata = 32'd17535;
			48002: outdata = 32'd17534;
			48003: outdata = 32'd17533;
			48004: outdata = 32'd17532;
			48005: outdata = 32'd17531;
			48006: outdata = 32'd17530;
			48007: outdata = 32'd17529;
			48008: outdata = 32'd17528;
			48009: outdata = 32'd17527;
			48010: outdata = 32'd17526;
			48011: outdata = 32'd17525;
			48012: outdata = 32'd17524;
			48013: outdata = 32'd17523;
			48014: outdata = 32'd17522;
			48015: outdata = 32'd17521;
			48016: outdata = 32'd17520;
			48017: outdata = 32'd17519;
			48018: outdata = 32'd17518;
			48019: outdata = 32'd17517;
			48020: outdata = 32'd17516;
			48021: outdata = 32'd17515;
			48022: outdata = 32'd17514;
			48023: outdata = 32'd17513;
			48024: outdata = 32'd17512;
			48025: outdata = 32'd17511;
			48026: outdata = 32'd17510;
			48027: outdata = 32'd17509;
			48028: outdata = 32'd17508;
			48029: outdata = 32'd17507;
			48030: outdata = 32'd17506;
			48031: outdata = 32'd17505;
			48032: outdata = 32'd17504;
			48033: outdata = 32'd17503;
			48034: outdata = 32'd17502;
			48035: outdata = 32'd17501;
			48036: outdata = 32'd17500;
			48037: outdata = 32'd17499;
			48038: outdata = 32'd17498;
			48039: outdata = 32'd17497;
			48040: outdata = 32'd17496;
			48041: outdata = 32'd17495;
			48042: outdata = 32'd17494;
			48043: outdata = 32'd17493;
			48044: outdata = 32'd17492;
			48045: outdata = 32'd17491;
			48046: outdata = 32'd17490;
			48047: outdata = 32'd17489;
			48048: outdata = 32'd17488;
			48049: outdata = 32'd17487;
			48050: outdata = 32'd17486;
			48051: outdata = 32'd17485;
			48052: outdata = 32'd17484;
			48053: outdata = 32'd17483;
			48054: outdata = 32'd17482;
			48055: outdata = 32'd17481;
			48056: outdata = 32'd17480;
			48057: outdata = 32'd17479;
			48058: outdata = 32'd17478;
			48059: outdata = 32'd17477;
			48060: outdata = 32'd17476;
			48061: outdata = 32'd17475;
			48062: outdata = 32'd17474;
			48063: outdata = 32'd17473;
			48064: outdata = 32'd17472;
			48065: outdata = 32'd17471;
			48066: outdata = 32'd17470;
			48067: outdata = 32'd17469;
			48068: outdata = 32'd17468;
			48069: outdata = 32'd17467;
			48070: outdata = 32'd17466;
			48071: outdata = 32'd17465;
			48072: outdata = 32'd17464;
			48073: outdata = 32'd17463;
			48074: outdata = 32'd17462;
			48075: outdata = 32'd17461;
			48076: outdata = 32'd17460;
			48077: outdata = 32'd17459;
			48078: outdata = 32'd17458;
			48079: outdata = 32'd17457;
			48080: outdata = 32'd17456;
			48081: outdata = 32'd17455;
			48082: outdata = 32'd17454;
			48083: outdata = 32'd17453;
			48084: outdata = 32'd17452;
			48085: outdata = 32'd17451;
			48086: outdata = 32'd17450;
			48087: outdata = 32'd17449;
			48088: outdata = 32'd17448;
			48089: outdata = 32'd17447;
			48090: outdata = 32'd17446;
			48091: outdata = 32'd17445;
			48092: outdata = 32'd17444;
			48093: outdata = 32'd17443;
			48094: outdata = 32'd17442;
			48095: outdata = 32'd17441;
			48096: outdata = 32'd17440;
			48097: outdata = 32'd17439;
			48098: outdata = 32'd17438;
			48099: outdata = 32'd17437;
			48100: outdata = 32'd17436;
			48101: outdata = 32'd17435;
			48102: outdata = 32'd17434;
			48103: outdata = 32'd17433;
			48104: outdata = 32'd17432;
			48105: outdata = 32'd17431;
			48106: outdata = 32'd17430;
			48107: outdata = 32'd17429;
			48108: outdata = 32'd17428;
			48109: outdata = 32'd17427;
			48110: outdata = 32'd17426;
			48111: outdata = 32'd17425;
			48112: outdata = 32'd17424;
			48113: outdata = 32'd17423;
			48114: outdata = 32'd17422;
			48115: outdata = 32'd17421;
			48116: outdata = 32'd17420;
			48117: outdata = 32'd17419;
			48118: outdata = 32'd17418;
			48119: outdata = 32'd17417;
			48120: outdata = 32'd17416;
			48121: outdata = 32'd17415;
			48122: outdata = 32'd17414;
			48123: outdata = 32'd17413;
			48124: outdata = 32'd17412;
			48125: outdata = 32'd17411;
			48126: outdata = 32'd17410;
			48127: outdata = 32'd17409;
			48128: outdata = 32'd17408;
			48129: outdata = 32'd17407;
			48130: outdata = 32'd17406;
			48131: outdata = 32'd17405;
			48132: outdata = 32'd17404;
			48133: outdata = 32'd17403;
			48134: outdata = 32'd17402;
			48135: outdata = 32'd17401;
			48136: outdata = 32'd17400;
			48137: outdata = 32'd17399;
			48138: outdata = 32'd17398;
			48139: outdata = 32'd17397;
			48140: outdata = 32'd17396;
			48141: outdata = 32'd17395;
			48142: outdata = 32'd17394;
			48143: outdata = 32'd17393;
			48144: outdata = 32'd17392;
			48145: outdata = 32'd17391;
			48146: outdata = 32'd17390;
			48147: outdata = 32'd17389;
			48148: outdata = 32'd17388;
			48149: outdata = 32'd17387;
			48150: outdata = 32'd17386;
			48151: outdata = 32'd17385;
			48152: outdata = 32'd17384;
			48153: outdata = 32'd17383;
			48154: outdata = 32'd17382;
			48155: outdata = 32'd17381;
			48156: outdata = 32'd17380;
			48157: outdata = 32'd17379;
			48158: outdata = 32'd17378;
			48159: outdata = 32'd17377;
			48160: outdata = 32'd17376;
			48161: outdata = 32'd17375;
			48162: outdata = 32'd17374;
			48163: outdata = 32'd17373;
			48164: outdata = 32'd17372;
			48165: outdata = 32'd17371;
			48166: outdata = 32'd17370;
			48167: outdata = 32'd17369;
			48168: outdata = 32'd17368;
			48169: outdata = 32'd17367;
			48170: outdata = 32'd17366;
			48171: outdata = 32'd17365;
			48172: outdata = 32'd17364;
			48173: outdata = 32'd17363;
			48174: outdata = 32'd17362;
			48175: outdata = 32'd17361;
			48176: outdata = 32'd17360;
			48177: outdata = 32'd17359;
			48178: outdata = 32'd17358;
			48179: outdata = 32'd17357;
			48180: outdata = 32'd17356;
			48181: outdata = 32'd17355;
			48182: outdata = 32'd17354;
			48183: outdata = 32'd17353;
			48184: outdata = 32'd17352;
			48185: outdata = 32'd17351;
			48186: outdata = 32'd17350;
			48187: outdata = 32'd17349;
			48188: outdata = 32'd17348;
			48189: outdata = 32'd17347;
			48190: outdata = 32'd17346;
			48191: outdata = 32'd17345;
			48192: outdata = 32'd17344;
			48193: outdata = 32'd17343;
			48194: outdata = 32'd17342;
			48195: outdata = 32'd17341;
			48196: outdata = 32'd17340;
			48197: outdata = 32'd17339;
			48198: outdata = 32'd17338;
			48199: outdata = 32'd17337;
			48200: outdata = 32'd17336;
			48201: outdata = 32'd17335;
			48202: outdata = 32'd17334;
			48203: outdata = 32'd17333;
			48204: outdata = 32'd17332;
			48205: outdata = 32'd17331;
			48206: outdata = 32'd17330;
			48207: outdata = 32'd17329;
			48208: outdata = 32'd17328;
			48209: outdata = 32'd17327;
			48210: outdata = 32'd17326;
			48211: outdata = 32'd17325;
			48212: outdata = 32'd17324;
			48213: outdata = 32'd17323;
			48214: outdata = 32'd17322;
			48215: outdata = 32'd17321;
			48216: outdata = 32'd17320;
			48217: outdata = 32'd17319;
			48218: outdata = 32'd17318;
			48219: outdata = 32'd17317;
			48220: outdata = 32'd17316;
			48221: outdata = 32'd17315;
			48222: outdata = 32'd17314;
			48223: outdata = 32'd17313;
			48224: outdata = 32'd17312;
			48225: outdata = 32'd17311;
			48226: outdata = 32'd17310;
			48227: outdata = 32'd17309;
			48228: outdata = 32'd17308;
			48229: outdata = 32'd17307;
			48230: outdata = 32'd17306;
			48231: outdata = 32'd17305;
			48232: outdata = 32'd17304;
			48233: outdata = 32'd17303;
			48234: outdata = 32'd17302;
			48235: outdata = 32'd17301;
			48236: outdata = 32'd17300;
			48237: outdata = 32'd17299;
			48238: outdata = 32'd17298;
			48239: outdata = 32'd17297;
			48240: outdata = 32'd17296;
			48241: outdata = 32'd17295;
			48242: outdata = 32'd17294;
			48243: outdata = 32'd17293;
			48244: outdata = 32'd17292;
			48245: outdata = 32'd17291;
			48246: outdata = 32'd17290;
			48247: outdata = 32'd17289;
			48248: outdata = 32'd17288;
			48249: outdata = 32'd17287;
			48250: outdata = 32'd17286;
			48251: outdata = 32'd17285;
			48252: outdata = 32'd17284;
			48253: outdata = 32'd17283;
			48254: outdata = 32'd17282;
			48255: outdata = 32'd17281;
			48256: outdata = 32'd17280;
			48257: outdata = 32'd17279;
			48258: outdata = 32'd17278;
			48259: outdata = 32'd17277;
			48260: outdata = 32'd17276;
			48261: outdata = 32'd17275;
			48262: outdata = 32'd17274;
			48263: outdata = 32'd17273;
			48264: outdata = 32'd17272;
			48265: outdata = 32'd17271;
			48266: outdata = 32'd17270;
			48267: outdata = 32'd17269;
			48268: outdata = 32'd17268;
			48269: outdata = 32'd17267;
			48270: outdata = 32'd17266;
			48271: outdata = 32'd17265;
			48272: outdata = 32'd17264;
			48273: outdata = 32'd17263;
			48274: outdata = 32'd17262;
			48275: outdata = 32'd17261;
			48276: outdata = 32'd17260;
			48277: outdata = 32'd17259;
			48278: outdata = 32'd17258;
			48279: outdata = 32'd17257;
			48280: outdata = 32'd17256;
			48281: outdata = 32'd17255;
			48282: outdata = 32'd17254;
			48283: outdata = 32'd17253;
			48284: outdata = 32'd17252;
			48285: outdata = 32'd17251;
			48286: outdata = 32'd17250;
			48287: outdata = 32'd17249;
			48288: outdata = 32'd17248;
			48289: outdata = 32'd17247;
			48290: outdata = 32'd17246;
			48291: outdata = 32'd17245;
			48292: outdata = 32'd17244;
			48293: outdata = 32'd17243;
			48294: outdata = 32'd17242;
			48295: outdata = 32'd17241;
			48296: outdata = 32'd17240;
			48297: outdata = 32'd17239;
			48298: outdata = 32'd17238;
			48299: outdata = 32'd17237;
			48300: outdata = 32'd17236;
			48301: outdata = 32'd17235;
			48302: outdata = 32'd17234;
			48303: outdata = 32'd17233;
			48304: outdata = 32'd17232;
			48305: outdata = 32'd17231;
			48306: outdata = 32'd17230;
			48307: outdata = 32'd17229;
			48308: outdata = 32'd17228;
			48309: outdata = 32'd17227;
			48310: outdata = 32'd17226;
			48311: outdata = 32'd17225;
			48312: outdata = 32'd17224;
			48313: outdata = 32'd17223;
			48314: outdata = 32'd17222;
			48315: outdata = 32'd17221;
			48316: outdata = 32'd17220;
			48317: outdata = 32'd17219;
			48318: outdata = 32'd17218;
			48319: outdata = 32'd17217;
			48320: outdata = 32'd17216;
			48321: outdata = 32'd17215;
			48322: outdata = 32'd17214;
			48323: outdata = 32'd17213;
			48324: outdata = 32'd17212;
			48325: outdata = 32'd17211;
			48326: outdata = 32'd17210;
			48327: outdata = 32'd17209;
			48328: outdata = 32'd17208;
			48329: outdata = 32'd17207;
			48330: outdata = 32'd17206;
			48331: outdata = 32'd17205;
			48332: outdata = 32'd17204;
			48333: outdata = 32'd17203;
			48334: outdata = 32'd17202;
			48335: outdata = 32'd17201;
			48336: outdata = 32'd17200;
			48337: outdata = 32'd17199;
			48338: outdata = 32'd17198;
			48339: outdata = 32'd17197;
			48340: outdata = 32'd17196;
			48341: outdata = 32'd17195;
			48342: outdata = 32'd17194;
			48343: outdata = 32'd17193;
			48344: outdata = 32'd17192;
			48345: outdata = 32'd17191;
			48346: outdata = 32'd17190;
			48347: outdata = 32'd17189;
			48348: outdata = 32'd17188;
			48349: outdata = 32'd17187;
			48350: outdata = 32'd17186;
			48351: outdata = 32'd17185;
			48352: outdata = 32'd17184;
			48353: outdata = 32'd17183;
			48354: outdata = 32'd17182;
			48355: outdata = 32'd17181;
			48356: outdata = 32'd17180;
			48357: outdata = 32'd17179;
			48358: outdata = 32'd17178;
			48359: outdata = 32'd17177;
			48360: outdata = 32'd17176;
			48361: outdata = 32'd17175;
			48362: outdata = 32'd17174;
			48363: outdata = 32'd17173;
			48364: outdata = 32'd17172;
			48365: outdata = 32'd17171;
			48366: outdata = 32'd17170;
			48367: outdata = 32'd17169;
			48368: outdata = 32'd17168;
			48369: outdata = 32'd17167;
			48370: outdata = 32'd17166;
			48371: outdata = 32'd17165;
			48372: outdata = 32'd17164;
			48373: outdata = 32'd17163;
			48374: outdata = 32'd17162;
			48375: outdata = 32'd17161;
			48376: outdata = 32'd17160;
			48377: outdata = 32'd17159;
			48378: outdata = 32'd17158;
			48379: outdata = 32'd17157;
			48380: outdata = 32'd17156;
			48381: outdata = 32'd17155;
			48382: outdata = 32'd17154;
			48383: outdata = 32'd17153;
			48384: outdata = 32'd17152;
			48385: outdata = 32'd17151;
			48386: outdata = 32'd17150;
			48387: outdata = 32'd17149;
			48388: outdata = 32'd17148;
			48389: outdata = 32'd17147;
			48390: outdata = 32'd17146;
			48391: outdata = 32'd17145;
			48392: outdata = 32'd17144;
			48393: outdata = 32'd17143;
			48394: outdata = 32'd17142;
			48395: outdata = 32'd17141;
			48396: outdata = 32'd17140;
			48397: outdata = 32'd17139;
			48398: outdata = 32'd17138;
			48399: outdata = 32'd17137;
			48400: outdata = 32'd17136;
			48401: outdata = 32'd17135;
			48402: outdata = 32'd17134;
			48403: outdata = 32'd17133;
			48404: outdata = 32'd17132;
			48405: outdata = 32'd17131;
			48406: outdata = 32'd17130;
			48407: outdata = 32'd17129;
			48408: outdata = 32'd17128;
			48409: outdata = 32'd17127;
			48410: outdata = 32'd17126;
			48411: outdata = 32'd17125;
			48412: outdata = 32'd17124;
			48413: outdata = 32'd17123;
			48414: outdata = 32'd17122;
			48415: outdata = 32'd17121;
			48416: outdata = 32'd17120;
			48417: outdata = 32'd17119;
			48418: outdata = 32'd17118;
			48419: outdata = 32'd17117;
			48420: outdata = 32'd17116;
			48421: outdata = 32'd17115;
			48422: outdata = 32'd17114;
			48423: outdata = 32'd17113;
			48424: outdata = 32'd17112;
			48425: outdata = 32'd17111;
			48426: outdata = 32'd17110;
			48427: outdata = 32'd17109;
			48428: outdata = 32'd17108;
			48429: outdata = 32'd17107;
			48430: outdata = 32'd17106;
			48431: outdata = 32'd17105;
			48432: outdata = 32'd17104;
			48433: outdata = 32'd17103;
			48434: outdata = 32'd17102;
			48435: outdata = 32'd17101;
			48436: outdata = 32'd17100;
			48437: outdata = 32'd17099;
			48438: outdata = 32'd17098;
			48439: outdata = 32'd17097;
			48440: outdata = 32'd17096;
			48441: outdata = 32'd17095;
			48442: outdata = 32'd17094;
			48443: outdata = 32'd17093;
			48444: outdata = 32'd17092;
			48445: outdata = 32'd17091;
			48446: outdata = 32'd17090;
			48447: outdata = 32'd17089;
			48448: outdata = 32'd17088;
			48449: outdata = 32'd17087;
			48450: outdata = 32'd17086;
			48451: outdata = 32'd17085;
			48452: outdata = 32'd17084;
			48453: outdata = 32'd17083;
			48454: outdata = 32'd17082;
			48455: outdata = 32'd17081;
			48456: outdata = 32'd17080;
			48457: outdata = 32'd17079;
			48458: outdata = 32'd17078;
			48459: outdata = 32'd17077;
			48460: outdata = 32'd17076;
			48461: outdata = 32'd17075;
			48462: outdata = 32'd17074;
			48463: outdata = 32'd17073;
			48464: outdata = 32'd17072;
			48465: outdata = 32'd17071;
			48466: outdata = 32'd17070;
			48467: outdata = 32'd17069;
			48468: outdata = 32'd17068;
			48469: outdata = 32'd17067;
			48470: outdata = 32'd17066;
			48471: outdata = 32'd17065;
			48472: outdata = 32'd17064;
			48473: outdata = 32'd17063;
			48474: outdata = 32'd17062;
			48475: outdata = 32'd17061;
			48476: outdata = 32'd17060;
			48477: outdata = 32'd17059;
			48478: outdata = 32'd17058;
			48479: outdata = 32'd17057;
			48480: outdata = 32'd17056;
			48481: outdata = 32'd17055;
			48482: outdata = 32'd17054;
			48483: outdata = 32'd17053;
			48484: outdata = 32'd17052;
			48485: outdata = 32'd17051;
			48486: outdata = 32'd17050;
			48487: outdata = 32'd17049;
			48488: outdata = 32'd17048;
			48489: outdata = 32'd17047;
			48490: outdata = 32'd17046;
			48491: outdata = 32'd17045;
			48492: outdata = 32'd17044;
			48493: outdata = 32'd17043;
			48494: outdata = 32'd17042;
			48495: outdata = 32'd17041;
			48496: outdata = 32'd17040;
			48497: outdata = 32'd17039;
			48498: outdata = 32'd17038;
			48499: outdata = 32'd17037;
			48500: outdata = 32'd17036;
			48501: outdata = 32'd17035;
			48502: outdata = 32'd17034;
			48503: outdata = 32'd17033;
			48504: outdata = 32'd17032;
			48505: outdata = 32'd17031;
			48506: outdata = 32'd17030;
			48507: outdata = 32'd17029;
			48508: outdata = 32'd17028;
			48509: outdata = 32'd17027;
			48510: outdata = 32'd17026;
			48511: outdata = 32'd17025;
			48512: outdata = 32'd17024;
			48513: outdata = 32'd17023;
			48514: outdata = 32'd17022;
			48515: outdata = 32'd17021;
			48516: outdata = 32'd17020;
			48517: outdata = 32'd17019;
			48518: outdata = 32'd17018;
			48519: outdata = 32'd17017;
			48520: outdata = 32'd17016;
			48521: outdata = 32'd17015;
			48522: outdata = 32'd17014;
			48523: outdata = 32'd17013;
			48524: outdata = 32'd17012;
			48525: outdata = 32'd17011;
			48526: outdata = 32'd17010;
			48527: outdata = 32'd17009;
			48528: outdata = 32'd17008;
			48529: outdata = 32'd17007;
			48530: outdata = 32'd17006;
			48531: outdata = 32'd17005;
			48532: outdata = 32'd17004;
			48533: outdata = 32'd17003;
			48534: outdata = 32'd17002;
			48535: outdata = 32'd17001;
			48536: outdata = 32'd17000;
			48537: outdata = 32'd16999;
			48538: outdata = 32'd16998;
			48539: outdata = 32'd16997;
			48540: outdata = 32'd16996;
			48541: outdata = 32'd16995;
			48542: outdata = 32'd16994;
			48543: outdata = 32'd16993;
			48544: outdata = 32'd16992;
			48545: outdata = 32'd16991;
			48546: outdata = 32'd16990;
			48547: outdata = 32'd16989;
			48548: outdata = 32'd16988;
			48549: outdata = 32'd16987;
			48550: outdata = 32'd16986;
			48551: outdata = 32'd16985;
			48552: outdata = 32'd16984;
			48553: outdata = 32'd16983;
			48554: outdata = 32'd16982;
			48555: outdata = 32'd16981;
			48556: outdata = 32'd16980;
			48557: outdata = 32'd16979;
			48558: outdata = 32'd16978;
			48559: outdata = 32'd16977;
			48560: outdata = 32'd16976;
			48561: outdata = 32'd16975;
			48562: outdata = 32'd16974;
			48563: outdata = 32'd16973;
			48564: outdata = 32'd16972;
			48565: outdata = 32'd16971;
			48566: outdata = 32'd16970;
			48567: outdata = 32'd16969;
			48568: outdata = 32'd16968;
			48569: outdata = 32'd16967;
			48570: outdata = 32'd16966;
			48571: outdata = 32'd16965;
			48572: outdata = 32'd16964;
			48573: outdata = 32'd16963;
			48574: outdata = 32'd16962;
			48575: outdata = 32'd16961;
			48576: outdata = 32'd16960;
			48577: outdata = 32'd16959;
			48578: outdata = 32'd16958;
			48579: outdata = 32'd16957;
			48580: outdata = 32'd16956;
			48581: outdata = 32'd16955;
			48582: outdata = 32'd16954;
			48583: outdata = 32'd16953;
			48584: outdata = 32'd16952;
			48585: outdata = 32'd16951;
			48586: outdata = 32'd16950;
			48587: outdata = 32'd16949;
			48588: outdata = 32'd16948;
			48589: outdata = 32'd16947;
			48590: outdata = 32'd16946;
			48591: outdata = 32'd16945;
			48592: outdata = 32'd16944;
			48593: outdata = 32'd16943;
			48594: outdata = 32'd16942;
			48595: outdata = 32'd16941;
			48596: outdata = 32'd16940;
			48597: outdata = 32'd16939;
			48598: outdata = 32'd16938;
			48599: outdata = 32'd16937;
			48600: outdata = 32'd16936;
			48601: outdata = 32'd16935;
			48602: outdata = 32'd16934;
			48603: outdata = 32'd16933;
			48604: outdata = 32'd16932;
			48605: outdata = 32'd16931;
			48606: outdata = 32'd16930;
			48607: outdata = 32'd16929;
			48608: outdata = 32'd16928;
			48609: outdata = 32'd16927;
			48610: outdata = 32'd16926;
			48611: outdata = 32'd16925;
			48612: outdata = 32'd16924;
			48613: outdata = 32'd16923;
			48614: outdata = 32'd16922;
			48615: outdata = 32'd16921;
			48616: outdata = 32'd16920;
			48617: outdata = 32'd16919;
			48618: outdata = 32'd16918;
			48619: outdata = 32'd16917;
			48620: outdata = 32'd16916;
			48621: outdata = 32'd16915;
			48622: outdata = 32'd16914;
			48623: outdata = 32'd16913;
			48624: outdata = 32'd16912;
			48625: outdata = 32'd16911;
			48626: outdata = 32'd16910;
			48627: outdata = 32'd16909;
			48628: outdata = 32'd16908;
			48629: outdata = 32'd16907;
			48630: outdata = 32'd16906;
			48631: outdata = 32'd16905;
			48632: outdata = 32'd16904;
			48633: outdata = 32'd16903;
			48634: outdata = 32'd16902;
			48635: outdata = 32'd16901;
			48636: outdata = 32'd16900;
			48637: outdata = 32'd16899;
			48638: outdata = 32'd16898;
			48639: outdata = 32'd16897;
			48640: outdata = 32'd16896;
			48641: outdata = 32'd16895;
			48642: outdata = 32'd16894;
			48643: outdata = 32'd16893;
			48644: outdata = 32'd16892;
			48645: outdata = 32'd16891;
			48646: outdata = 32'd16890;
			48647: outdata = 32'd16889;
			48648: outdata = 32'd16888;
			48649: outdata = 32'd16887;
			48650: outdata = 32'd16886;
			48651: outdata = 32'd16885;
			48652: outdata = 32'd16884;
			48653: outdata = 32'd16883;
			48654: outdata = 32'd16882;
			48655: outdata = 32'd16881;
			48656: outdata = 32'd16880;
			48657: outdata = 32'd16879;
			48658: outdata = 32'd16878;
			48659: outdata = 32'd16877;
			48660: outdata = 32'd16876;
			48661: outdata = 32'd16875;
			48662: outdata = 32'd16874;
			48663: outdata = 32'd16873;
			48664: outdata = 32'd16872;
			48665: outdata = 32'd16871;
			48666: outdata = 32'd16870;
			48667: outdata = 32'd16869;
			48668: outdata = 32'd16868;
			48669: outdata = 32'd16867;
			48670: outdata = 32'd16866;
			48671: outdata = 32'd16865;
			48672: outdata = 32'd16864;
			48673: outdata = 32'd16863;
			48674: outdata = 32'd16862;
			48675: outdata = 32'd16861;
			48676: outdata = 32'd16860;
			48677: outdata = 32'd16859;
			48678: outdata = 32'd16858;
			48679: outdata = 32'd16857;
			48680: outdata = 32'd16856;
			48681: outdata = 32'd16855;
			48682: outdata = 32'd16854;
			48683: outdata = 32'd16853;
			48684: outdata = 32'd16852;
			48685: outdata = 32'd16851;
			48686: outdata = 32'd16850;
			48687: outdata = 32'd16849;
			48688: outdata = 32'd16848;
			48689: outdata = 32'd16847;
			48690: outdata = 32'd16846;
			48691: outdata = 32'd16845;
			48692: outdata = 32'd16844;
			48693: outdata = 32'd16843;
			48694: outdata = 32'd16842;
			48695: outdata = 32'd16841;
			48696: outdata = 32'd16840;
			48697: outdata = 32'd16839;
			48698: outdata = 32'd16838;
			48699: outdata = 32'd16837;
			48700: outdata = 32'd16836;
			48701: outdata = 32'd16835;
			48702: outdata = 32'd16834;
			48703: outdata = 32'd16833;
			48704: outdata = 32'd16832;
			48705: outdata = 32'd16831;
			48706: outdata = 32'd16830;
			48707: outdata = 32'd16829;
			48708: outdata = 32'd16828;
			48709: outdata = 32'd16827;
			48710: outdata = 32'd16826;
			48711: outdata = 32'd16825;
			48712: outdata = 32'd16824;
			48713: outdata = 32'd16823;
			48714: outdata = 32'd16822;
			48715: outdata = 32'd16821;
			48716: outdata = 32'd16820;
			48717: outdata = 32'd16819;
			48718: outdata = 32'd16818;
			48719: outdata = 32'd16817;
			48720: outdata = 32'd16816;
			48721: outdata = 32'd16815;
			48722: outdata = 32'd16814;
			48723: outdata = 32'd16813;
			48724: outdata = 32'd16812;
			48725: outdata = 32'd16811;
			48726: outdata = 32'd16810;
			48727: outdata = 32'd16809;
			48728: outdata = 32'd16808;
			48729: outdata = 32'd16807;
			48730: outdata = 32'd16806;
			48731: outdata = 32'd16805;
			48732: outdata = 32'd16804;
			48733: outdata = 32'd16803;
			48734: outdata = 32'd16802;
			48735: outdata = 32'd16801;
			48736: outdata = 32'd16800;
			48737: outdata = 32'd16799;
			48738: outdata = 32'd16798;
			48739: outdata = 32'd16797;
			48740: outdata = 32'd16796;
			48741: outdata = 32'd16795;
			48742: outdata = 32'd16794;
			48743: outdata = 32'd16793;
			48744: outdata = 32'd16792;
			48745: outdata = 32'd16791;
			48746: outdata = 32'd16790;
			48747: outdata = 32'd16789;
			48748: outdata = 32'd16788;
			48749: outdata = 32'd16787;
			48750: outdata = 32'd16786;
			48751: outdata = 32'd16785;
			48752: outdata = 32'd16784;
			48753: outdata = 32'd16783;
			48754: outdata = 32'd16782;
			48755: outdata = 32'd16781;
			48756: outdata = 32'd16780;
			48757: outdata = 32'd16779;
			48758: outdata = 32'd16778;
			48759: outdata = 32'd16777;
			48760: outdata = 32'd16776;
			48761: outdata = 32'd16775;
			48762: outdata = 32'd16774;
			48763: outdata = 32'd16773;
			48764: outdata = 32'd16772;
			48765: outdata = 32'd16771;
			48766: outdata = 32'd16770;
			48767: outdata = 32'd16769;
			48768: outdata = 32'd16768;
			48769: outdata = 32'd16767;
			48770: outdata = 32'd16766;
			48771: outdata = 32'd16765;
			48772: outdata = 32'd16764;
			48773: outdata = 32'd16763;
			48774: outdata = 32'd16762;
			48775: outdata = 32'd16761;
			48776: outdata = 32'd16760;
			48777: outdata = 32'd16759;
			48778: outdata = 32'd16758;
			48779: outdata = 32'd16757;
			48780: outdata = 32'd16756;
			48781: outdata = 32'd16755;
			48782: outdata = 32'd16754;
			48783: outdata = 32'd16753;
			48784: outdata = 32'd16752;
			48785: outdata = 32'd16751;
			48786: outdata = 32'd16750;
			48787: outdata = 32'd16749;
			48788: outdata = 32'd16748;
			48789: outdata = 32'd16747;
			48790: outdata = 32'd16746;
			48791: outdata = 32'd16745;
			48792: outdata = 32'd16744;
			48793: outdata = 32'd16743;
			48794: outdata = 32'd16742;
			48795: outdata = 32'd16741;
			48796: outdata = 32'd16740;
			48797: outdata = 32'd16739;
			48798: outdata = 32'd16738;
			48799: outdata = 32'd16737;
			48800: outdata = 32'd16736;
			48801: outdata = 32'd16735;
			48802: outdata = 32'd16734;
			48803: outdata = 32'd16733;
			48804: outdata = 32'd16732;
			48805: outdata = 32'd16731;
			48806: outdata = 32'd16730;
			48807: outdata = 32'd16729;
			48808: outdata = 32'd16728;
			48809: outdata = 32'd16727;
			48810: outdata = 32'd16726;
			48811: outdata = 32'd16725;
			48812: outdata = 32'd16724;
			48813: outdata = 32'd16723;
			48814: outdata = 32'd16722;
			48815: outdata = 32'd16721;
			48816: outdata = 32'd16720;
			48817: outdata = 32'd16719;
			48818: outdata = 32'd16718;
			48819: outdata = 32'd16717;
			48820: outdata = 32'd16716;
			48821: outdata = 32'd16715;
			48822: outdata = 32'd16714;
			48823: outdata = 32'd16713;
			48824: outdata = 32'd16712;
			48825: outdata = 32'd16711;
			48826: outdata = 32'd16710;
			48827: outdata = 32'd16709;
			48828: outdata = 32'd16708;
			48829: outdata = 32'd16707;
			48830: outdata = 32'd16706;
			48831: outdata = 32'd16705;
			48832: outdata = 32'd16704;
			48833: outdata = 32'd16703;
			48834: outdata = 32'd16702;
			48835: outdata = 32'd16701;
			48836: outdata = 32'd16700;
			48837: outdata = 32'd16699;
			48838: outdata = 32'd16698;
			48839: outdata = 32'd16697;
			48840: outdata = 32'd16696;
			48841: outdata = 32'd16695;
			48842: outdata = 32'd16694;
			48843: outdata = 32'd16693;
			48844: outdata = 32'd16692;
			48845: outdata = 32'd16691;
			48846: outdata = 32'd16690;
			48847: outdata = 32'd16689;
			48848: outdata = 32'd16688;
			48849: outdata = 32'd16687;
			48850: outdata = 32'd16686;
			48851: outdata = 32'd16685;
			48852: outdata = 32'd16684;
			48853: outdata = 32'd16683;
			48854: outdata = 32'd16682;
			48855: outdata = 32'd16681;
			48856: outdata = 32'd16680;
			48857: outdata = 32'd16679;
			48858: outdata = 32'd16678;
			48859: outdata = 32'd16677;
			48860: outdata = 32'd16676;
			48861: outdata = 32'd16675;
			48862: outdata = 32'd16674;
			48863: outdata = 32'd16673;
			48864: outdata = 32'd16672;
			48865: outdata = 32'd16671;
			48866: outdata = 32'd16670;
			48867: outdata = 32'd16669;
			48868: outdata = 32'd16668;
			48869: outdata = 32'd16667;
			48870: outdata = 32'd16666;
			48871: outdata = 32'd16665;
			48872: outdata = 32'd16664;
			48873: outdata = 32'd16663;
			48874: outdata = 32'd16662;
			48875: outdata = 32'd16661;
			48876: outdata = 32'd16660;
			48877: outdata = 32'd16659;
			48878: outdata = 32'd16658;
			48879: outdata = 32'd16657;
			48880: outdata = 32'd16656;
			48881: outdata = 32'd16655;
			48882: outdata = 32'd16654;
			48883: outdata = 32'd16653;
			48884: outdata = 32'd16652;
			48885: outdata = 32'd16651;
			48886: outdata = 32'd16650;
			48887: outdata = 32'd16649;
			48888: outdata = 32'd16648;
			48889: outdata = 32'd16647;
			48890: outdata = 32'd16646;
			48891: outdata = 32'd16645;
			48892: outdata = 32'd16644;
			48893: outdata = 32'd16643;
			48894: outdata = 32'd16642;
			48895: outdata = 32'd16641;
			48896: outdata = 32'd16640;
			48897: outdata = 32'd16639;
			48898: outdata = 32'd16638;
			48899: outdata = 32'd16637;
			48900: outdata = 32'd16636;
			48901: outdata = 32'd16635;
			48902: outdata = 32'd16634;
			48903: outdata = 32'd16633;
			48904: outdata = 32'd16632;
			48905: outdata = 32'd16631;
			48906: outdata = 32'd16630;
			48907: outdata = 32'd16629;
			48908: outdata = 32'd16628;
			48909: outdata = 32'd16627;
			48910: outdata = 32'd16626;
			48911: outdata = 32'd16625;
			48912: outdata = 32'd16624;
			48913: outdata = 32'd16623;
			48914: outdata = 32'd16622;
			48915: outdata = 32'd16621;
			48916: outdata = 32'd16620;
			48917: outdata = 32'd16619;
			48918: outdata = 32'd16618;
			48919: outdata = 32'd16617;
			48920: outdata = 32'd16616;
			48921: outdata = 32'd16615;
			48922: outdata = 32'd16614;
			48923: outdata = 32'd16613;
			48924: outdata = 32'd16612;
			48925: outdata = 32'd16611;
			48926: outdata = 32'd16610;
			48927: outdata = 32'd16609;
			48928: outdata = 32'd16608;
			48929: outdata = 32'd16607;
			48930: outdata = 32'd16606;
			48931: outdata = 32'd16605;
			48932: outdata = 32'd16604;
			48933: outdata = 32'd16603;
			48934: outdata = 32'd16602;
			48935: outdata = 32'd16601;
			48936: outdata = 32'd16600;
			48937: outdata = 32'd16599;
			48938: outdata = 32'd16598;
			48939: outdata = 32'd16597;
			48940: outdata = 32'd16596;
			48941: outdata = 32'd16595;
			48942: outdata = 32'd16594;
			48943: outdata = 32'd16593;
			48944: outdata = 32'd16592;
			48945: outdata = 32'd16591;
			48946: outdata = 32'd16590;
			48947: outdata = 32'd16589;
			48948: outdata = 32'd16588;
			48949: outdata = 32'd16587;
			48950: outdata = 32'd16586;
			48951: outdata = 32'd16585;
			48952: outdata = 32'd16584;
			48953: outdata = 32'd16583;
			48954: outdata = 32'd16582;
			48955: outdata = 32'd16581;
			48956: outdata = 32'd16580;
			48957: outdata = 32'd16579;
			48958: outdata = 32'd16578;
			48959: outdata = 32'd16577;
			48960: outdata = 32'd16576;
			48961: outdata = 32'd16575;
			48962: outdata = 32'd16574;
			48963: outdata = 32'd16573;
			48964: outdata = 32'd16572;
			48965: outdata = 32'd16571;
			48966: outdata = 32'd16570;
			48967: outdata = 32'd16569;
			48968: outdata = 32'd16568;
			48969: outdata = 32'd16567;
			48970: outdata = 32'd16566;
			48971: outdata = 32'd16565;
			48972: outdata = 32'd16564;
			48973: outdata = 32'd16563;
			48974: outdata = 32'd16562;
			48975: outdata = 32'd16561;
			48976: outdata = 32'd16560;
			48977: outdata = 32'd16559;
			48978: outdata = 32'd16558;
			48979: outdata = 32'd16557;
			48980: outdata = 32'd16556;
			48981: outdata = 32'd16555;
			48982: outdata = 32'd16554;
			48983: outdata = 32'd16553;
			48984: outdata = 32'd16552;
			48985: outdata = 32'd16551;
			48986: outdata = 32'd16550;
			48987: outdata = 32'd16549;
			48988: outdata = 32'd16548;
			48989: outdata = 32'd16547;
			48990: outdata = 32'd16546;
			48991: outdata = 32'd16545;
			48992: outdata = 32'd16544;
			48993: outdata = 32'd16543;
			48994: outdata = 32'd16542;
			48995: outdata = 32'd16541;
			48996: outdata = 32'd16540;
			48997: outdata = 32'd16539;
			48998: outdata = 32'd16538;
			48999: outdata = 32'd16537;
			49000: outdata = 32'd16536;
			49001: outdata = 32'd16535;
			49002: outdata = 32'd16534;
			49003: outdata = 32'd16533;
			49004: outdata = 32'd16532;
			49005: outdata = 32'd16531;
			49006: outdata = 32'd16530;
			49007: outdata = 32'd16529;
			49008: outdata = 32'd16528;
			49009: outdata = 32'd16527;
			49010: outdata = 32'd16526;
			49011: outdata = 32'd16525;
			49012: outdata = 32'd16524;
			49013: outdata = 32'd16523;
			49014: outdata = 32'd16522;
			49015: outdata = 32'd16521;
			49016: outdata = 32'd16520;
			49017: outdata = 32'd16519;
			49018: outdata = 32'd16518;
			49019: outdata = 32'd16517;
			49020: outdata = 32'd16516;
			49021: outdata = 32'd16515;
			49022: outdata = 32'd16514;
			49023: outdata = 32'd16513;
			49024: outdata = 32'd16512;
			49025: outdata = 32'd16511;
			49026: outdata = 32'd16510;
			49027: outdata = 32'd16509;
			49028: outdata = 32'd16508;
			49029: outdata = 32'd16507;
			49030: outdata = 32'd16506;
			49031: outdata = 32'd16505;
			49032: outdata = 32'd16504;
			49033: outdata = 32'd16503;
			49034: outdata = 32'd16502;
			49035: outdata = 32'd16501;
			49036: outdata = 32'd16500;
			49037: outdata = 32'd16499;
			49038: outdata = 32'd16498;
			49039: outdata = 32'd16497;
			49040: outdata = 32'd16496;
			49041: outdata = 32'd16495;
			49042: outdata = 32'd16494;
			49043: outdata = 32'd16493;
			49044: outdata = 32'd16492;
			49045: outdata = 32'd16491;
			49046: outdata = 32'd16490;
			49047: outdata = 32'd16489;
			49048: outdata = 32'd16488;
			49049: outdata = 32'd16487;
			49050: outdata = 32'd16486;
			49051: outdata = 32'd16485;
			49052: outdata = 32'd16484;
			49053: outdata = 32'd16483;
			49054: outdata = 32'd16482;
			49055: outdata = 32'd16481;
			49056: outdata = 32'd16480;
			49057: outdata = 32'd16479;
			49058: outdata = 32'd16478;
			49059: outdata = 32'd16477;
			49060: outdata = 32'd16476;
			49061: outdata = 32'd16475;
			49062: outdata = 32'd16474;
			49063: outdata = 32'd16473;
			49064: outdata = 32'd16472;
			49065: outdata = 32'd16471;
			49066: outdata = 32'd16470;
			49067: outdata = 32'd16469;
			49068: outdata = 32'd16468;
			49069: outdata = 32'd16467;
			49070: outdata = 32'd16466;
			49071: outdata = 32'd16465;
			49072: outdata = 32'd16464;
			49073: outdata = 32'd16463;
			49074: outdata = 32'd16462;
			49075: outdata = 32'd16461;
			49076: outdata = 32'd16460;
			49077: outdata = 32'd16459;
			49078: outdata = 32'd16458;
			49079: outdata = 32'd16457;
			49080: outdata = 32'd16456;
			49081: outdata = 32'd16455;
			49082: outdata = 32'd16454;
			49083: outdata = 32'd16453;
			49084: outdata = 32'd16452;
			49085: outdata = 32'd16451;
			49086: outdata = 32'd16450;
			49087: outdata = 32'd16449;
			49088: outdata = 32'd16448;
			49089: outdata = 32'd16447;
			49090: outdata = 32'd16446;
			49091: outdata = 32'd16445;
			49092: outdata = 32'd16444;
			49093: outdata = 32'd16443;
			49094: outdata = 32'd16442;
			49095: outdata = 32'd16441;
			49096: outdata = 32'd16440;
			49097: outdata = 32'd16439;
			49098: outdata = 32'd16438;
			49099: outdata = 32'd16437;
			49100: outdata = 32'd16436;
			49101: outdata = 32'd16435;
			49102: outdata = 32'd16434;
			49103: outdata = 32'd16433;
			49104: outdata = 32'd16432;
			49105: outdata = 32'd16431;
			49106: outdata = 32'd16430;
			49107: outdata = 32'd16429;
			49108: outdata = 32'd16428;
			49109: outdata = 32'd16427;
			49110: outdata = 32'd16426;
			49111: outdata = 32'd16425;
			49112: outdata = 32'd16424;
			49113: outdata = 32'd16423;
			49114: outdata = 32'd16422;
			49115: outdata = 32'd16421;
			49116: outdata = 32'd16420;
			49117: outdata = 32'd16419;
			49118: outdata = 32'd16418;
			49119: outdata = 32'd16417;
			49120: outdata = 32'd16416;
			49121: outdata = 32'd16415;
			49122: outdata = 32'd16414;
			49123: outdata = 32'd16413;
			49124: outdata = 32'd16412;
			49125: outdata = 32'd16411;
			49126: outdata = 32'd16410;
			49127: outdata = 32'd16409;
			49128: outdata = 32'd16408;
			49129: outdata = 32'd16407;
			49130: outdata = 32'd16406;
			49131: outdata = 32'd16405;
			49132: outdata = 32'd16404;
			49133: outdata = 32'd16403;
			49134: outdata = 32'd16402;
			49135: outdata = 32'd16401;
			49136: outdata = 32'd16400;
			49137: outdata = 32'd16399;
			49138: outdata = 32'd16398;
			49139: outdata = 32'd16397;
			49140: outdata = 32'd16396;
			49141: outdata = 32'd16395;
			49142: outdata = 32'd16394;
			49143: outdata = 32'd16393;
			49144: outdata = 32'd16392;
			49145: outdata = 32'd16391;
			49146: outdata = 32'd16390;
			49147: outdata = 32'd16389;
			49148: outdata = 32'd16388;
			49149: outdata = 32'd16387;
			49150: outdata = 32'd16386;
			49151: outdata = 32'd16385;
			49152: outdata = 32'd16384;
			49153: outdata = 32'd16383;
			49154: outdata = 32'd16382;
			49155: outdata = 32'd16381;
			49156: outdata = 32'd16380;
			49157: outdata = 32'd16379;
			49158: outdata = 32'd16378;
			49159: outdata = 32'd16377;
			49160: outdata = 32'd16376;
			49161: outdata = 32'd16375;
			49162: outdata = 32'd16374;
			49163: outdata = 32'd16373;
			49164: outdata = 32'd16372;
			49165: outdata = 32'd16371;
			49166: outdata = 32'd16370;
			49167: outdata = 32'd16369;
			49168: outdata = 32'd16368;
			49169: outdata = 32'd16367;
			49170: outdata = 32'd16366;
			49171: outdata = 32'd16365;
			49172: outdata = 32'd16364;
			49173: outdata = 32'd16363;
			49174: outdata = 32'd16362;
			49175: outdata = 32'd16361;
			49176: outdata = 32'd16360;
			49177: outdata = 32'd16359;
			49178: outdata = 32'd16358;
			49179: outdata = 32'd16357;
			49180: outdata = 32'd16356;
			49181: outdata = 32'd16355;
			49182: outdata = 32'd16354;
			49183: outdata = 32'd16353;
			49184: outdata = 32'd16352;
			49185: outdata = 32'd16351;
			49186: outdata = 32'd16350;
			49187: outdata = 32'd16349;
			49188: outdata = 32'd16348;
			49189: outdata = 32'd16347;
			49190: outdata = 32'd16346;
			49191: outdata = 32'd16345;
			49192: outdata = 32'd16344;
			49193: outdata = 32'd16343;
			49194: outdata = 32'd16342;
			49195: outdata = 32'd16341;
			49196: outdata = 32'd16340;
			49197: outdata = 32'd16339;
			49198: outdata = 32'd16338;
			49199: outdata = 32'd16337;
			49200: outdata = 32'd16336;
			49201: outdata = 32'd16335;
			49202: outdata = 32'd16334;
			49203: outdata = 32'd16333;
			49204: outdata = 32'd16332;
			49205: outdata = 32'd16331;
			49206: outdata = 32'd16330;
			49207: outdata = 32'd16329;
			49208: outdata = 32'd16328;
			49209: outdata = 32'd16327;
			49210: outdata = 32'd16326;
			49211: outdata = 32'd16325;
			49212: outdata = 32'd16324;
			49213: outdata = 32'd16323;
			49214: outdata = 32'd16322;
			49215: outdata = 32'd16321;
			49216: outdata = 32'd16320;
			49217: outdata = 32'd16319;
			49218: outdata = 32'd16318;
			49219: outdata = 32'd16317;
			49220: outdata = 32'd16316;
			49221: outdata = 32'd16315;
			49222: outdata = 32'd16314;
			49223: outdata = 32'd16313;
			49224: outdata = 32'd16312;
			49225: outdata = 32'd16311;
			49226: outdata = 32'd16310;
			49227: outdata = 32'd16309;
			49228: outdata = 32'd16308;
			49229: outdata = 32'd16307;
			49230: outdata = 32'd16306;
			49231: outdata = 32'd16305;
			49232: outdata = 32'd16304;
			49233: outdata = 32'd16303;
			49234: outdata = 32'd16302;
			49235: outdata = 32'd16301;
			49236: outdata = 32'd16300;
			49237: outdata = 32'd16299;
			49238: outdata = 32'd16298;
			49239: outdata = 32'd16297;
			49240: outdata = 32'd16296;
			49241: outdata = 32'd16295;
			49242: outdata = 32'd16294;
			49243: outdata = 32'd16293;
			49244: outdata = 32'd16292;
			49245: outdata = 32'd16291;
			49246: outdata = 32'd16290;
			49247: outdata = 32'd16289;
			49248: outdata = 32'd16288;
			49249: outdata = 32'd16287;
			49250: outdata = 32'd16286;
			49251: outdata = 32'd16285;
			49252: outdata = 32'd16284;
			49253: outdata = 32'd16283;
			49254: outdata = 32'd16282;
			49255: outdata = 32'd16281;
			49256: outdata = 32'd16280;
			49257: outdata = 32'd16279;
			49258: outdata = 32'd16278;
			49259: outdata = 32'd16277;
			49260: outdata = 32'd16276;
			49261: outdata = 32'd16275;
			49262: outdata = 32'd16274;
			49263: outdata = 32'd16273;
			49264: outdata = 32'd16272;
			49265: outdata = 32'd16271;
			49266: outdata = 32'd16270;
			49267: outdata = 32'd16269;
			49268: outdata = 32'd16268;
			49269: outdata = 32'd16267;
			49270: outdata = 32'd16266;
			49271: outdata = 32'd16265;
			49272: outdata = 32'd16264;
			49273: outdata = 32'd16263;
			49274: outdata = 32'd16262;
			49275: outdata = 32'd16261;
			49276: outdata = 32'd16260;
			49277: outdata = 32'd16259;
			49278: outdata = 32'd16258;
			49279: outdata = 32'd16257;
			49280: outdata = 32'd16256;
			49281: outdata = 32'd16255;
			49282: outdata = 32'd16254;
			49283: outdata = 32'd16253;
			49284: outdata = 32'd16252;
			49285: outdata = 32'd16251;
			49286: outdata = 32'd16250;
			49287: outdata = 32'd16249;
			49288: outdata = 32'd16248;
			49289: outdata = 32'd16247;
			49290: outdata = 32'd16246;
			49291: outdata = 32'd16245;
			49292: outdata = 32'd16244;
			49293: outdata = 32'd16243;
			49294: outdata = 32'd16242;
			49295: outdata = 32'd16241;
			49296: outdata = 32'd16240;
			49297: outdata = 32'd16239;
			49298: outdata = 32'd16238;
			49299: outdata = 32'd16237;
			49300: outdata = 32'd16236;
			49301: outdata = 32'd16235;
			49302: outdata = 32'd16234;
			49303: outdata = 32'd16233;
			49304: outdata = 32'd16232;
			49305: outdata = 32'd16231;
			49306: outdata = 32'd16230;
			49307: outdata = 32'd16229;
			49308: outdata = 32'd16228;
			49309: outdata = 32'd16227;
			49310: outdata = 32'd16226;
			49311: outdata = 32'd16225;
			49312: outdata = 32'd16224;
			49313: outdata = 32'd16223;
			49314: outdata = 32'd16222;
			49315: outdata = 32'd16221;
			49316: outdata = 32'd16220;
			49317: outdata = 32'd16219;
			49318: outdata = 32'd16218;
			49319: outdata = 32'd16217;
			49320: outdata = 32'd16216;
			49321: outdata = 32'd16215;
			49322: outdata = 32'd16214;
			49323: outdata = 32'd16213;
			49324: outdata = 32'd16212;
			49325: outdata = 32'd16211;
			49326: outdata = 32'd16210;
			49327: outdata = 32'd16209;
			49328: outdata = 32'd16208;
			49329: outdata = 32'd16207;
			49330: outdata = 32'd16206;
			49331: outdata = 32'd16205;
			49332: outdata = 32'd16204;
			49333: outdata = 32'd16203;
			49334: outdata = 32'd16202;
			49335: outdata = 32'd16201;
			49336: outdata = 32'd16200;
			49337: outdata = 32'd16199;
			49338: outdata = 32'd16198;
			49339: outdata = 32'd16197;
			49340: outdata = 32'd16196;
			49341: outdata = 32'd16195;
			49342: outdata = 32'd16194;
			49343: outdata = 32'd16193;
			49344: outdata = 32'd16192;
			49345: outdata = 32'd16191;
			49346: outdata = 32'd16190;
			49347: outdata = 32'd16189;
			49348: outdata = 32'd16188;
			49349: outdata = 32'd16187;
			49350: outdata = 32'd16186;
			49351: outdata = 32'd16185;
			49352: outdata = 32'd16184;
			49353: outdata = 32'd16183;
			49354: outdata = 32'd16182;
			49355: outdata = 32'd16181;
			49356: outdata = 32'd16180;
			49357: outdata = 32'd16179;
			49358: outdata = 32'd16178;
			49359: outdata = 32'd16177;
			49360: outdata = 32'd16176;
			49361: outdata = 32'd16175;
			49362: outdata = 32'd16174;
			49363: outdata = 32'd16173;
			49364: outdata = 32'd16172;
			49365: outdata = 32'd16171;
			49366: outdata = 32'd16170;
			49367: outdata = 32'd16169;
			49368: outdata = 32'd16168;
			49369: outdata = 32'd16167;
			49370: outdata = 32'd16166;
			49371: outdata = 32'd16165;
			49372: outdata = 32'd16164;
			49373: outdata = 32'd16163;
			49374: outdata = 32'd16162;
			49375: outdata = 32'd16161;
			49376: outdata = 32'd16160;
			49377: outdata = 32'd16159;
			49378: outdata = 32'd16158;
			49379: outdata = 32'd16157;
			49380: outdata = 32'd16156;
			49381: outdata = 32'd16155;
			49382: outdata = 32'd16154;
			49383: outdata = 32'd16153;
			49384: outdata = 32'd16152;
			49385: outdata = 32'd16151;
			49386: outdata = 32'd16150;
			49387: outdata = 32'd16149;
			49388: outdata = 32'd16148;
			49389: outdata = 32'd16147;
			49390: outdata = 32'd16146;
			49391: outdata = 32'd16145;
			49392: outdata = 32'd16144;
			49393: outdata = 32'd16143;
			49394: outdata = 32'd16142;
			49395: outdata = 32'd16141;
			49396: outdata = 32'd16140;
			49397: outdata = 32'd16139;
			49398: outdata = 32'd16138;
			49399: outdata = 32'd16137;
			49400: outdata = 32'd16136;
			49401: outdata = 32'd16135;
			49402: outdata = 32'd16134;
			49403: outdata = 32'd16133;
			49404: outdata = 32'd16132;
			49405: outdata = 32'd16131;
			49406: outdata = 32'd16130;
			49407: outdata = 32'd16129;
			49408: outdata = 32'd16128;
			49409: outdata = 32'd16127;
			49410: outdata = 32'd16126;
			49411: outdata = 32'd16125;
			49412: outdata = 32'd16124;
			49413: outdata = 32'd16123;
			49414: outdata = 32'd16122;
			49415: outdata = 32'd16121;
			49416: outdata = 32'd16120;
			49417: outdata = 32'd16119;
			49418: outdata = 32'd16118;
			49419: outdata = 32'd16117;
			49420: outdata = 32'd16116;
			49421: outdata = 32'd16115;
			49422: outdata = 32'd16114;
			49423: outdata = 32'd16113;
			49424: outdata = 32'd16112;
			49425: outdata = 32'd16111;
			49426: outdata = 32'd16110;
			49427: outdata = 32'd16109;
			49428: outdata = 32'd16108;
			49429: outdata = 32'd16107;
			49430: outdata = 32'd16106;
			49431: outdata = 32'd16105;
			49432: outdata = 32'd16104;
			49433: outdata = 32'd16103;
			49434: outdata = 32'd16102;
			49435: outdata = 32'd16101;
			49436: outdata = 32'd16100;
			49437: outdata = 32'd16099;
			49438: outdata = 32'd16098;
			49439: outdata = 32'd16097;
			49440: outdata = 32'd16096;
			49441: outdata = 32'd16095;
			49442: outdata = 32'd16094;
			49443: outdata = 32'd16093;
			49444: outdata = 32'd16092;
			49445: outdata = 32'd16091;
			49446: outdata = 32'd16090;
			49447: outdata = 32'd16089;
			49448: outdata = 32'd16088;
			49449: outdata = 32'd16087;
			49450: outdata = 32'd16086;
			49451: outdata = 32'd16085;
			49452: outdata = 32'd16084;
			49453: outdata = 32'd16083;
			49454: outdata = 32'd16082;
			49455: outdata = 32'd16081;
			49456: outdata = 32'd16080;
			49457: outdata = 32'd16079;
			49458: outdata = 32'd16078;
			49459: outdata = 32'd16077;
			49460: outdata = 32'd16076;
			49461: outdata = 32'd16075;
			49462: outdata = 32'd16074;
			49463: outdata = 32'd16073;
			49464: outdata = 32'd16072;
			49465: outdata = 32'd16071;
			49466: outdata = 32'd16070;
			49467: outdata = 32'd16069;
			49468: outdata = 32'd16068;
			49469: outdata = 32'd16067;
			49470: outdata = 32'd16066;
			49471: outdata = 32'd16065;
			49472: outdata = 32'd16064;
			49473: outdata = 32'd16063;
			49474: outdata = 32'd16062;
			49475: outdata = 32'd16061;
			49476: outdata = 32'd16060;
			49477: outdata = 32'd16059;
			49478: outdata = 32'd16058;
			49479: outdata = 32'd16057;
			49480: outdata = 32'd16056;
			49481: outdata = 32'd16055;
			49482: outdata = 32'd16054;
			49483: outdata = 32'd16053;
			49484: outdata = 32'd16052;
			49485: outdata = 32'd16051;
			49486: outdata = 32'd16050;
			49487: outdata = 32'd16049;
			49488: outdata = 32'd16048;
			49489: outdata = 32'd16047;
			49490: outdata = 32'd16046;
			49491: outdata = 32'd16045;
			49492: outdata = 32'd16044;
			49493: outdata = 32'd16043;
			49494: outdata = 32'd16042;
			49495: outdata = 32'd16041;
			49496: outdata = 32'd16040;
			49497: outdata = 32'd16039;
			49498: outdata = 32'd16038;
			49499: outdata = 32'd16037;
			49500: outdata = 32'd16036;
			49501: outdata = 32'd16035;
			49502: outdata = 32'd16034;
			49503: outdata = 32'd16033;
			49504: outdata = 32'd16032;
			49505: outdata = 32'd16031;
			49506: outdata = 32'd16030;
			49507: outdata = 32'd16029;
			49508: outdata = 32'd16028;
			49509: outdata = 32'd16027;
			49510: outdata = 32'd16026;
			49511: outdata = 32'd16025;
			49512: outdata = 32'd16024;
			49513: outdata = 32'd16023;
			49514: outdata = 32'd16022;
			49515: outdata = 32'd16021;
			49516: outdata = 32'd16020;
			49517: outdata = 32'd16019;
			49518: outdata = 32'd16018;
			49519: outdata = 32'd16017;
			49520: outdata = 32'd16016;
			49521: outdata = 32'd16015;
			49522: outdata = 32'd16014;
			49523: outdata = 32'd16013;
			49524: outdata = 32'd16012;
			49525: outdata = 32'd16011;
			49526: outdata = 32'd16010;
			49527: outdata = 32'd16009;
			49528: outdata = 32'd16008;
			49529: outdata = 32'd16007;
			49530: outdata = 32'd16006;
			49531: outdata = 32'd16005;
			49532: outdata = 32'd16004;
			49533: outdata = 32'd16003;
			49534: outdata = 32'd16002;
			49535: outdata = 32'd16001;
			49536: outdata = 32'd16000;
			49537: outdata = 32'd15999;
			49538: outdata = 32'd15998;
			49539: outdata = 32'd15997;
			49540: outdata = 32'd15996;
			49541: outdata = 32'd15995;
			49542: outdata = 32'd15994;
			49543: outdata = 32'd15993;
			49544: outdata = 32'd15992;
			49545: outdata = 32'd15991;
			49546: outdata = 32'd15990;
			49547: outdata = 32'd15989;
			49548: outdata = 32'd15988;
			49549: outdata = 32'd15987;
			49550: outdata = 32'd15986;
			49551: outdata = 32'd15985;
			49552: outdata = 32'd15984;
			49553: outdata = 32'd15983;
			49554: outdata = 32'd15982;
			49555: outdata = 32'd15981;
			49556: outdata = 32'd15980;
			49557: outdata = 32'd15979;
			49558: outdata = 32'd15978;
			49559: outdata = 32'd15977;
			49560: outdata = 32'd15976;
			49561: outdata = 32'd15975;
			49562: outdata = 32'd15974;
			49563: outdata = 32'd15973;
			49564: outdata = 32'd15972;
			49565: outdata = 32'd15971;
			49566: outdata = 32'd15970;
			49567: outdata = 32'd15969;
			49568: outdata = 32'd15968;
			49569: outdata = 32'd15967;
			49570: outdata = 32'd15966;
			49571: outdata = 32'd15965;
			49572: outdata = 32'd15964;
			49573: outdata = 32'd15963;
			49574: outdata = 32'd15962;
			49575: outdata = 32'd15961;
			49576: outdata = 32'd15960;
			49577: outdata = 32'd15959;
			49578: outdata = 32'd15958;
			49579: outdata = 32'd15957;
			49580: outdata = 32'd15956;
			49581: outdata = 32'd15955;
			49582: outdata = 32'd15954;
			49583: outdata = 32'd15953;
			49584: outdata = 32'd15952;
			49585: outdata = 32'd15951;
			49586: outdata = 32'd15950;
			49587: outdata = 32'd15949;
			49588: outdata = 32'd15948;
			49589: outdata = 32'd15947;
			49590: outdata = 32'd15946;
			49591: outdata = 32'd15945;
			49592: outdata = 32'd15944;
			49593: outdata = 32'd15943;
			49594: outdata = 32'd15942;
			49595: outdata = 32'd15941;
			49596: outdata = 32'd15940;
			49597: outdata = 32'd15939;
			49598: outdata = 32'd15938;
			49599: outdata = 32'd15937;
			49600: outdata = 32'd15936;
			49601: outdata = 32'd15935;
			49602: outdata = 32'd15934;
			49603: outdata = 32'd15933;
			49604: outdata = 32'd15932;
			49605: outdata = 32'd15931;
			49606: outdata = 32'd15930;
			49607: outdata = 32'd15929;
			49608: outdata = 32'd15928;
			49609: outdata = 32'd15927;
			49610: outdata = 32'd15926;
			49611: outdata = 32'd15925;
			49612: outdata = 32'd15924;
			49613: outdata = 32'd15923;
			49614: outdata = 32'd15922;
			49615: outdata = 32'd15921;
			49616: outdata = 32'd15920;
			49617: outdata = 32'd15919;
			49618: outdata = 32'd15918;
			49619: outdata = 32'd15917;
			49620: outdata = 32'd15916;
			49621: outdata = 32'd15915;
			49622: outdata = 32'd15914;
			49623: outdata = 32'd15913;
			49624: outdata = 32'd15912;
			49625: outdata = 32'd15911;
			49626: outdata = 32'd15910;
			49627: outdata = 32'd15909;
			49628: outdata = 32'd15908;
			49629: outdata = 32'd15907;
			49630: outdata = 32'd15906;
			49631: outdata = 32'd15905;
			49632: outdata = 32'd15904;
			49633: outdata = 32'd15903;
			49634: outdata = 32'd15902;
			49635: outdata = 32'd15901;
			49636: outdata = 32'd15900;
			49637: outdata = 32'd15899;
			49638: outdata = 32'd15898;
			49639: outdata = 32'd15897;
			49640: outdata = 32'd15896;
			49641: outdata = 32'd15895;
			49642: outdata = 32'd15894;
			49643: outdata = 32'd15893;
			49644: outdata = 32'd15892;
			49645: outdata = 32'd15891;
			49646: outdata = 32'd15890;
			49647: outdata = 32'd15889;
			49648: outdata = 32'd15888;
			49649: outdata = 32'd15887;
			49650: outdata = 32'd15886;
			49651: outdata = 32'd15885;
			49652: outdata = 32'd15884;
			49653: outdata = 32'd15883;
			49654: outdata = 32'd15882;
			49655: outdata = 32'd15881;
			49656: outdata = 32'd15880;
			49657: outdata = 32'd15879;
			49658: outdata = 32'd15878;
			49659: outdata = 32'd15877;
			49660: outdata = 32'd15876;
			49661: outdata = 32'd15875;
			49662: outdata = 32'd15874;
			49663: outdata = 32'd15873;
			49664: outdata = 32'd15872;
			49665: outdata = 32'd15871;
			49666: outdata = 32'd15870;
			49667: outdata = 32'd15869;
			49668: outdata = 32'd15868;
			49669: outdata = 32'd15867;
			49670: outdata = 32'd15866;
			49671: outdata = 32'd15865;
			49672: outdata = 32'd15864;
			49673: outdata = 32'd15863;
			49674: outdata = 32'd15862;
			49675: outdata = 32'd15861;
			49676: outdata = 32'd15860;
			49677: outdata = 32'd15859;
			49678: outdata = 32'd15858;
			49679: outdata = 32'd15857;
			49680: outdata = 32'd15856;
			49681: outdata = 32'd15855;
			49682: outdata = 32'd15854;
			49683: outdata = 32'd15853;
			49684: outdata = 32'd15852;
			49685: outdata = 32'd15851;
			49686: outdata = 32'd15850;
			49687: outdata = 32'd15849;
			49688: outdata = 32'd15848;
			49689: outdata = 32'd15847;
			49690: outdata = 32'd15846;
			49691: outdata = 32'd15845;
			49692: outdata = 32'd15844;
			49693: outdata = 32'd15843;
			49694: outdata = 32'd15842;
			49695: outdata = 32'd15841;
			49696: outdata = 32'd15840;
			49697: outdata = 32'd15839;
			49698: outdata = 32'd15838;
			49699: outdata = 32'd15837;
			49700: outdata = 32'd15836;
			49701: outdata = 32'd15835;
			49702: outdata = 32'd15834;
			49703: outdata = 32'd15833;
			49704: outdata = 32'd15832;
			49705: outdata = 32'd15831;
			49706: outdata = 32'd15830;
			49707: outdata = 32'd15829;
			49708: outdata = 32'd15828;
			49709: outdata = 32'd15827;
			49710: outdata = 32'd15826;
			49711: outdata = 32'd15825;
			49712: outdata = 32'd15824;
			49713: outdata = 32'd15823;
			49714: outdata = 32'd15822;
			49715: outdata = 32'd15821;
			49716: outdata = 32'd15820;
			49717: outdata = 32'd15819;
			49718: outdata = 32'd15818;
			49719: outdata = 32'd15817;
			49720: outdata = 32'd15816;
			49721: outdata = 32'd15815;
			49722: outdata = 32'd15814;
			49723: outdata = 32'd15813;
			49724: outdata = 32'd15812;
			49725: outdata = 32'd15811;
			49726: outdata = 32'd15810;
			49727: outdata = 32'd15809;
			49728: outdata = 32'd15808;
			49729: outdata = 32'd15807;
			49730: outdata = 32'd15806;
			49731: outdata = 32'd15805;
			49732: outdata = 32'd15804;
			49733: outdata = 32'd15803;
			49734: outdata = 32'd15802;
			49735: outdata = 32'd15801;
			49736: outdata = 32'd15800;
			49737: outdata = 32'd15799;
			49738: outdata = 32'd15798;
			49739: outdata = 32'd15797;
			49740: outdata = 32'd15796;
			49741: outdata = 32'd15795;
			49742: outdata = 32'd15794;
			49743: outdata = 32'd15793;
			49744: outdata = 32'd15792;
			49745: outdata = 32'd15791;
			49746: outdata = 32'd15790;
			49747: outdata = 32'd15789;
			49748: outdata = 32'd15788;
			49749: outdata = 32'd15787;
			49750: outdata = 32'd15786;
			49751: outdata = 32'd15785;
			49752: outdata = 32'd15784;
			49753: outdata = 32'd15783;
			49754: outdata = 32'd15782;
			49755: outdata = 32'd15781;
			49756: outdata = 32'd15780;
			49757: outdata = 32'd15779;
			49758: outdata = 32'd15778;
			49759: outdata = 32'd15777;
			49760: outdata = 32'd15776;
			49761: outdata = 32'd15775;
			49762: outdata = 32'd15774;
			49763: outdata = 32'd15773;
			49764: outdata = 32'd15772;
			49765: outdata = 32'd15771;
			49766: outdata = 32'd15770;
			49767: outdata = 32'd15769;
			49768: outdata = 32'd15768;
			49769: outdata = 32'd15767;
			49770: outdata = 32'd15766;
			49771: outdata = 32'd15765;
			49772: outdata = 32'd15764;
			49773: outdata = 32'd15763;
			49774: outdata = 32'd15762;
			49775: outdata = 32'd15761;
			49776: outdata = 32'd15760;
			49777: outdata = 32'd15759;
			49778: outdata = 32'd15758;
			49779: outdata = 32'd15757;
			49780: outdata = 32'd15756;
			49781: outdata = 32'd15755;
			49782: outdata = 32'd15754;
			49783: outdata = 32'd15753;
			49784: outdata = 32'd15752;
			49785: outdata = 32'd15751;
			49786: outdata = 32'd15750;
			49787: outdata = 32'd15749;
			49788: outdata = 32'd15748;
			49789: outdata = 32'd15747;
			49790: outdata = 32'd15746;
			49791: outdata = 32'd15745;
			49792: outdata = 32'd15744;
			49793: outdata = 32'd15743;
			49794: outdata = 32'd15742;
			49795: outdata = 32'd15741;
			49796: outdata = 32'd15740;
			49797: outdata = 32'd15739;
			49798: outdata = 32'd15738;
			49799: outdata = 32'd15737;
			49800: outdata = 32'd15736;
			49801: outdata = 32'd15735;
			49802: outdata = 32'd15734;
			49803: outdata = 32'd15733;
			49804: outdata = 32'd15732;
			49805: outdata = 32'd15731;
			49806: outdata = 32'd15730;
			49807: outdata = 32'd15729;
			49808: outdata = 32'd15728;
			49809: outdata = 32'd15727;
			49810: outdata = 32'd15726;
			49811: outdata = 32'd15725;
			49812: outdata = 32'd15724;
			49813: outdata = 32'd15723;
			49814: outdata = 32'd15722;
			49815: outdata = 32'd15721;
			49816: outdata = 32'd15720;
			49817: outdata = 32'd15719;
			49818: outdata = 32'd15718;
			49819: outdata = 32'd15717;
			49820: outdata = 32'd15716;
			49821: outdata = 32'd15715;
			49822: outdata = 32'd15714;
			49823: outdata = 32'd15713;
			49824: outdata = 32'd15712;
			49825: outdata = 32'd15711;
			49826: outdata = 32'd15710;
			49827: outdata = 32'd15709;
			49828: outdata = 32'd15708;
			49829: outdata = 32'd15707;
			49830: outdata = 32'd15706;
			49831: outdata = 32'd15705;
			49832: outdata = 32'd15704;
			49833: outdata = 32'd15703;
			49834: outdata = 32'd15702;
			49835: outdata = 32'd15701;
			49836: outdata = 32'd15700;
			49837: outdata = 32'd15699;
			49838: outdata = 32'd15698;
			49839: outdata = 32'd15697;
			49840: outdata = 32'd15696;
			49841: outdata = 32'd15695;
			49842: outdata = 32'd15694;
			49843: outdata = 32'd15693;
			49844: outdata = 32'd15692;
			49845: outdata = 32'd15691;
			49846: outdata = 32'd15690;
			49847: outdata = 32'd15689;
			49848: outdata = 32'd15688;
			49849: outdata = 32'd15687;
			49850: outdata = 32'd15686;
			49851: outdata = 32'd15685;
			49852: outdata = 32'd15684;
			49853: outdata = 32'd15683;
			49854: outdata = 32'd15682;
			49855: outdata = 32'd15681;
			49856: outdata = 32'd15680;
			49857: outdata = 32'd15679;
			49858: outdata = 32'd15678;
			49859: outdata = 32'd15677;
			49860: outdata = 32'd15676;
			49861: outdata = 32'd15675;
			49862: outdata = 32'd15674;
			49863: outdata = 32'd15673;
			49864: outdata = 32'd15672;
			49865: outdata = 32'd15671;
			49866: outdata = 32'd15670;
			49867: outdata = 32'd15669;
			49868: outdata = 32'd15668;
			49869: outdata = 32'd15667;
			49870: outdata = 32'd15666;
			49871: outdata = 32'd15665;
			49872: outdata = 32'd15664;
			49873: outdata = 32'd15663;
			49874: outdata = 32'd15662;
			49875: outdata = 32'd15661;
			49876: outdata = 32'd15660;
			49877: outdata = 32'd15659;
			49878: outdata = 32'd15658;
			49879: outdata = 32'd15657;
			49880: outdata = 32'd15656;
			49881: outdata = 32'd15655;
			49882: outdata = 32'd15654;
			49883: outdata = 32'd15653;
			49884: outdata = 32'd15652;
			49885: outdata = 32'd15651;
			49886: outdata = 32'd15650;
			49887: outdata = 32'd15649;
			49888: outdata = 32'd15648;
			49889: outdata = 32'd15647;
			49890: outdata = 32'd15646;
			49891: outdata = 32'd15645;
			49892: outdata = 32'd15644;
			49893: outdata = 32'd15643;
			49894: outdata = 32'd15642;
			49895: outdata = 32'd15641;
			49896: outdata = 32'd15640;
			49897: outdata = 32'd15639;
			49898: outdata = 32'd15638;
			49899: outdata = 32'd15637;
			49900: outdata = 32'd15636;
			49901: outdata = 32'd15635;
			49902: outdata = 32'd15634;
			49903: outdata = 32'd15633;
			49904: outdata = 32'd15632;
			49905: outdata = 32'd15631;
			49906: outdata = 32'd15630;
			49907: outdata = 32'd15629;
			49908: outdata = 32'd15628;
			49909: outdata = 32'd15627;
			49910: outdata = 32'd15626;
			49911: outdata = 32'd15625;
			49912: outdata = 32'd15624;
			49913: outdata = 32'd15623;
			49914: outdata = 32'd15622;
			49915: outdata = 32'd15621;
			49916: outdata = 32'd15620;
			49917: outdata = 32'd15619;
			49918: outdata = 32'd15618;
			49919: outdata = 32'd15617;
			49920: outdata = 32'd15616;
			49921: outdata = 32'd15615;
			49922: outdata = 32'd15614;
			49923: outdata = 32'd15613;
			49924: outdata = 32'd15612;
			49925: outdata = 32'd15611;
			49926: outdata = 32'd15610;
			49927: outdata = 32'd15609;
			49928: outdata = 32'd15608;
			49929: outdata = 32'd15607;
			49930: outdata = 32'd15606;
			49931: outdata = 32'd15605;
			49932: outdata = 32'd15604;
			49933: outdata = 32'd15603;
			49934: outdata = 32'd15602;
			49935: outdata = 32'd15601;
			49936: outdata = 32'd15600;
			49937: outdata = 32'd15599;
			49938: outdata = 32'd15598;
			49939: outdata = 32'd15597;
			49940: outdata = 32'd15596;
			49941: outdata = 32'd15595;
			49942: outdata = 32'd15594;
			49943: outdata = 32'd15593;
			49944: outdata = 32'd15592;
			49945: outdata = 32'd15591;
			49946: outdata = 32'd15590;
			49947: outdata = 32'd15589;
			49948: outdata = 32'd15588;
			49949: outdata = 32'd15587;
			49950: outdata = 32'd15586;
			49951: outdata = 32'd15585;
			49952: outdata = 32'd15584;
			49953: outdata = 32'd15583;
			49954: outdata = 32'd15582;
			49955: outdata = 32'd15581;
			49956: outdata = 32'd15580;
			49957: outdata = 32'd15579;
			49958: outdata = 32'd15578;
			49959: outdata = 32'd15577;
			49960: outdata = 32'd15576;
			49961: outdata = 32'd15575;
			49962: outdata = 32'd15574;
			49963: outdata = 32'd15573;
			49964: outdata = 32'd15572;
			49965: outdata = 32'd15571;
			49966: outdata = 32'd15570;
			49967: outdata = 32'd15569;
			49968: outdata = 32'd15568;
			49969: outdata = 32'd15567;
			49970: outdata = 32'd15566;
			49971: outdata = 32'd15565;
			49972: outdata = 32'd15564;
			49973: outdata = 32'd15563;
			49974: outdata = 32'd15562;
			49975: outdata = 32'd15561;
			49976: outdata = 32'd15560;
			49977: outdata = 32'd15559;
			49978: outdata = 32'd15558;
			49979: outdata = 32'd15557;
			49980: outdata = 32'd15556;
			49981: outdata = 32'd15555;
			49982: outdata = 32'd15554;
			49983: outdata = 32'd15553;
			49984: outdata = 32'd15552;
			49985: outdata = 32'd15551;
			49986: outdata = 32'd15550;
			49987: outdata = 32'd15549;
			49988: outdata = 32'd15548;
			49989: outdata = 32'd15547;
			49990: outdata = 32'd15546;
			49991: outdata = 32'd15545;
			49992: outdata = 32'd15544;
			49993: outdata = 32'd15543;
			49994: outdata = 32'd15542;
			49995: outdata = 32'd15541;
			49996: outdata = 32'd15540;
			49997: outdata = 32'd15539;
			49998: outdata = 32'd15538;
			49999: outdata = 32'd15537;
			50000: outdata = 32'd15536;
			50001: outdata = 32'd15535;
			50002: outdata = 32'd15534;
			50003: outdata = 32'd15533;
			50004: outdata = 32'd15532;
			50005: outdata = 32'd15531;
			50006: outdata = 32'd15530;
			50007: outdata = 32'd15529;
			50008: outdata = 32'd15528;
			50009: outdata = 32'd15527;
			50010: outdata = 32'd15526;
			50011: outdata = 32'd15525;
			50012: outdata = 32'd15524;
			50013: outdata = 32'd15523;
			50014: outdata = 32'd15522;
			50015: outdata = 32'd15521;
			50016: outdata = 32'd15520;
			50017: outdata = 32'd15519;
			50018: outdata = 32'd15518;
			50019: outdata = 32'd15517;
			50020: outdata = 32'd15516;
			50021: outdata = 32'd15515;
			50022: outdata = 32'd15514;
			50023: outdata = 32'd15513;
			50024: outdata = 32'd15512;
			50025: outdata = 32'd15511;
			50026: outdata = 32'd15510;
			50027: outdata = 32'd15509;
			50028: outdata = 32'd15508;
			50029: outdata = 32'd15507;
			50030: outdata = 32'd15506;
			50031: outdata = 32'd15505;
			50032: outdata = 32'd15504;
			50033: outdata = 32'd15503;
			50034: outdata = 32'd15502;
			50035: outdata = 32'd15501;
			50036: outdata = 32'd15500;
			50037: outdata = 32'd15499;
			50038: outdata = 32'd15498;
			50039: outdata = 32'd15497;
			50040: outdata = 32'd15496;
			50041: outdata = 32'd15495;
			50042: outdata = 32'd15494;
			50043: outdata = 32'd15493;
			50044: outdata = 32'd15492;
			50045: outdata = 32'd15491;
			50046: outdata = 32'd15490;
			50047: outdata = 32'd15489;
			50048: outdata = 32'd15488;
			50049: outdata = 32'd15487;
			50050: outdata = 32'd15486;
			50051: outdata = 32'd15485;
			50052: outdata = 32'd15484;
			50053: outdata = 32'd15483;
			50054: outdata = 32'd15482;
			50055: outdata = 32'd15481;
			50056: outdata = 32'd15480;
			50057: outdata = 32'd15479;
			50058: outdata = 32'd15478;
			50059: outdata = 32'd15477;
			50060: outdata = 32'd15476;
			50061: outdata = 32'd15475;
			50062: outdata = 32'd15474;
			50063: outdata = 32'd15473;
			50064: outdata = 32'd15472;
			50065: outdata = 32'd15471;
			50066: outdata = 32'd15470;
			50067: outdata = 32'd15469;
			50068: outdata = 32'd15468;
			50069: outdata = 32'd15467;
			50070: outdata = 32'd15466;
			50071: outdata = 32'd15465;
			50072: outdata = 32'd15464;
			50073: outdata = 32'd15463;
			50074: outdata = 32'd15462;
			50075: outdata = 32'd15461;
			50076: outdata = 32'd15460;
			50077: outdata = 32'd15459;
			50078: outdata = 32'd15458;
			50079: outdata = 32'd15457;
			50080: outdata = 32'd15456;
			50081: outdata = 32'd15455;
			50082: outdata = 32'd15454;
			50083: outdata = 32'd15453;
			50084: outdata = 32'd15452;
			50085: outdata = 32'd15451;
			50086: outdata = 32'd15450;
			50087: outdata = 32'd15449;
			50088: outdata = 32'd15448;
			50089: outdata = 32'd15447;
			50090: outdata = 32'd15446;
			50091: outdata = 32'd15445;
			50092: outdata = 32'd15444;
			50093: outdata = 32'd15443;
			50094: outdata = 32'd15442;
			50095: outdata = 32'd15441;
			50096: outdata = 32'd15440;
			50097: outdata = 32'd15439;
			50098: outdata = 32'd15438;
			50099: outdata = 32'd15437;
			50100: outdata = 32'd15436;
			50101: outdata = 32'd15435;
			50102: outdata = 32'd15434;
			50103: outdata = 32'd15433;
			50104: outdata = 32'd15432;
			50105: outdata = 32'd15431;
			50106: outdata = 32'd15430;
			50107: outdata = 32'd15429;
			50108: outdata = 32'd15428;
			50109: outdata = 32'd15427;
			50110: outdata = 32'd15426;
			50111: outdata = 32'd15425;
			50112: outdata = 32'd15424;
			50113: outdata = 32'd15423;
			50114: outdata = 32'd15422;
			50115: outdata = 32'd15421;
			50116: outdata = 32'd15420;
			50117: outdata = 32'd15419;
			50118: outdata = 32'd15418;
			50119: outdata = 32'd15417;
			50120: outdata = 32'd15416;
			50121: outdata = 32'd15415;
			50122: outdata = 32'd15414;
			50123: outdata = 32'd15413;
			50124: outdata = 32'd15412;
			50125: outdata = 32'd15411;
			50126: outdata = 32'd15410;
			50127: outdata = 32'd15409;
			50128: outdata = 32'd15408;
			50129: outdata = 32'd15407;
			50130: outdata = 32'd15406;
			50131: outdata = 32'd15405;
			50132: outdata = 32'd15404;
			50133: outdata = 32'd15403;
			50134: outdata = 32'd15402;
			50135: outdata = 32'd15401;
			50136: outdata = 32'd15400;
			50137: outdata = 32'd15399;
			50138: outdata = 32'd15398;
			50139: outdata = 32'd15397;
			50140: outdata = 32'd15396;
			50141: outdata = 32'd15395;
			50142: outdata = 32'd15394;
			50143: outdata = 32'd15393;
			50144: outdata = 32'd15392;
			50145: outdata = 32'd15391;
			50146: outdata = 32'd15390;
			50147: outdata = 32'd15389;
			50148: outdata = 32'd15388;
			50149: outdata = 32'd15387;
			50150: outdata = 32'd15386;
			50151: outdata = 32'd15385;
			50152: outdata = 32'd15384;
			50153: outdata = 32'd15383;
			50154: outdata = 32'd15382;
			50155: outdata = 32'd15381;
			50156: outdata = 32'd15380;
			50157: outdata = 32'd15379;
			50158: outdata = 32'd15378;
			50159: outdata = 32'd15377;
			50160: outdata = 32'd15376;
			50161: outdata = 32'd15375;
			50162: outdata = 32'd15374;
			50163: outdata = 32'd15373;
			50164: outdata = 32'd15372;
			50165: outdata = 32'd15371;
			50166: outdata = 32'd15370;
			50167: outdata = 32'd15369;
			50168: outdata = 32'd15368;
			50169: outdata = 32'd15367;
			50170: outdata = 32'd15366;
			50171: outdata = 32'd15365;
			50172: outdata = 32'd15364;
			50173: outdata = 32'd15363;
			50174: outdata = 32'd15362;
			50175: outdata = 32'd15361;
			50176: outdata = 32'd15360;
			50177: outdata = 32'd15359;
			50178: outdata = 32'd15358;
			50179: outdata = 32'd15357;
			50180: outdata = 32'd15356;
			50181: outdata = 32'd15355;
			50182: outdata = 32'd15354;
			50183: outdata = 32'd15353;
			50184: outdata = 32'd15352;
			50185: outdata = 32'd15351;
			50186: outdata = 32'd15350;
			50187: outdata = 32'd15349;
			50188: outdata = 32'd15348;
			50189: outdata = 32'd15347;
			50190: outdata = 32'd15346;
			50191: outdata = 32'd15345;
			50192: outdata = 32'd15344;
			50193: outdata = 32'd15343;
			50194: outdata = 32'd15342;
			50195: outdata = 32'd15341;
			50196: outdata = 32'd15340;
			50197: outdata = 32'd15339;
			50198: outdata = 32'd15338;
			50199: outdata = 32'd15337;
			50200: outdata = 32'd15336;
			50201: outdata = 32'd15335;
			50202: outdata = 32'd15334;
			50203: outdata = 32'd15333;
			50204: outdata = 32'd15332;
			50205: outdata = 32'd15331;
			50206: outdata = 32'd15330;
			50207: outdata = 32'd15329;
			50208: outdata = 32'd15328;
			50209: outdata = 32'd15327;
			50210: outdata = 32'd15326;
			50211: outdata = 32'd15325;
			50212: outdata = 32'd15324;
			50213: outdata = 32'd15323;
			50214: outdata = 32'd15322;
			50215: outdata = 32'd15321;
			50216: outdata = 32'd15320;
			50217: outdata = 32'd15319;
			50218: outdata = 32'd15318;
			50219: outdata = 32'd15317;
			50220: outdata = 32'd15316;
			50221: outdata = 32'd15315;
			50222: outdata = 32'd15314;
			50223: outdata = 32'd15313;
			50224: outdata = 32'd15312;
			50225: outdata = 32'd15311;
			50226: outdata = 32'd15310;
			50227: outdata = 32'd15309;
			50228: outdata = 32'd15308;
			50229: outdata = 32'd15307;
			50230: outdata = 32'd15306;
			50231: outdata = 32'd15305;
			50232: outdata = 32'd15304;
			50233: outdata = 32'd15303;
			50234: outdata = 32'd15302;
			50235: outdata = 32'd15301;
			50236: outdata = 32'd15300;
			50237: outdata = 32'd15299;
			50238: outdata = 32'd15298;
			50239: outdata = 32'd15297;
			50240: outdata = 32'd15296;
			50241: outdata = 32'd15295;
			50242: outdata = 32'd15294;
			50243: outdata = 32'd15293;
			50244: outdata = 32'd15292;
			50245: outdata = 32'd15291;
			50246: outdata = 32'd15290;
			50247: outdata = 32'd15289;
			50248: outdata = 32'd15288;
			50249: outdata = 32'd15287;
			50250: outdata = 32'd15286;
			50251: outdata = 32'd15285;
			50252: outdata = 32'd15284;
			50253: outdata = 32'd15283;
			50254: outdata = 32'd15282;
			50255: outdata = 32'd15281;
			50256: outdata = 32'd15280;
			50257: outdata = 32'd15279;
			50258: outdata = 32'd15278;
			50259: outdata = 32'd15277;
			50260: outdata = 32'd15276;
			50261: outdata = 32'd15275;
			50262: outdata = 32'd15274;
			50263: outdata = 32'd15273;
			50264: outdata = 32'd15272;
			50265: outdata = 32'd15271;
			50266: outdata = 32'd15270;
			50267: outdata = 32'd15269;
			50268: outdata = 32'd15268;
			50269: outdata = 32'd15267;
			50270: outdata = 32'd15266;
			50271: outdata = 32'd15265;
			50272: outdata = 32'd15264;
			50273: outdata = 32'd15263;
			50274: outdata = 32'd15262;
			50275: outdata = 32'd15261;
			50276: outdata = 32'd15260;
			50277: outdata = 32'd15259;
			50278: outdata = 32'd15258;
			50279: outdata = 32'd15257;
			50280: outdata = 32'd15256;
			50281: outdata = 32'd15255;
			50282: outdata = 32'd15254;
			50283: outdata = 32'd15253;
			50284: outdata = 32'd15252;
			50285: outdata = 32'd15251;
			50286: outdata = 32'd15250;
			50287: outdata = 32'd15249;
			50288: outdata = 32'd15248;
			50289: outdata = 32'd15247;
			50290: outdata = 32'd15246;
			50291: outdata = 32'd15245;
			50292: outdata = 32'd15244;
			50293: outdata = 32'd15243;
			50294: outdata = 32'd15242;
			50295: outdata = 32'd15241;
			50296: outdata = 32'd15240;
			50297: outdata = 32'd15239;
			50298: outdata = 32'd15238;
			50299: outdata = 32'd15237;
			50300: outdata = 32'd15236;
			50301: outdata = 32'd15235;
			50302: outdata = 32'd15234;
			50303: outdata = 32'd15233;
			50304: outdata = 32'd15232;
			50305: outdata = 32'd15231;
			50306: outdata = 32'd15230;
			50307: outdata = 32'd15229;
			50308: outdata = 32'd15228;
			50309: outdata = 32'd15227;
			50310: outdata = 32'd15226;
			50311: outdata = 32'd15225;
			50312: outdata = 32'd15224;
			50313: outdata = 32'd15223;
			50314: outdata = 32'd15222;
			50315: outdata = 32'd15221;
			50316: outdata = 32'd15220;
			50317: outdata = 32'd15219;
			50318: outdata = 32'd15218;
			50319: outdata = 32'd15217;
			50320: outdata = 32'd15216;
			50321: outdata = 32'd15215;
			50322: outdata = 32'd15214;
			50323: outdata = 32'd15213;
			50324: outdata = 32'd15212;
			50325: outdata = 32'd15211;
			50326: outdata = 32'd15210;
			50327: outdata = 32'd15209;
			50328: outdata = 32'd15208;
			50329: outdata = 32'd15207;
			50330: outdata = 32'd15206;
			50331: outdata = 32'd15205;
			50332: outdata = 32'd15204;
			50333: outdata = 32'd15203;
			50334: outdata = 32'd15202;
			50335: outdata = 32'd15201;
			50336: outdata = 32'd15200;
			50337: outdata = 32'd15199;
			50338: outdata = 32'd15198;
			50339: outdata = 32'd15197;
			50340: outdata = 32'd15196;
			50341: outdata = 32'd15195;
			50342: outdata = 32'd15194;
			50343: outdata = 32'd15193;
			50344: outdata = 32'd15192;
			50345: outdata = 32'd15191;
			50346: outdata = 32'd15190;
			50347: outdata = 32'd15189;
			50348: outdata = 32'd15188;
			50349: outdata = 32'd15187;
			50350: outdata = 32'd15186;
			50351: outdata = 32'd15185;
			50352: outdata = 32'd15184;
			50353: outdata = 32'd15183;
			50354: outdata = 32'd15182;
			50355: outdata = 32'd15181;
			50356: outdata = 32'd15180;
			50357: outdata = 32'd15179;
			50358: outdata = 32'd15178;
			50359: outdata = 32'd15177;
			50360: outdata = 32'd15176;
			50361: outdata = 32'd15175;
			50362: outdata = 32'd15174;
			50363: outdata = 32'd15173;
			50364: outdata = 32'd15172;
			50365: outdata = 32'd15171;
			50366: outdata = 32'd15170;
			50367: outdata = 32'd15169;
			50368: outdata = 32'd15168;
			50369: outdata = 32'd15167;
			50370: outdata = 32'd15166;
			50371: outdata = 32'd15165;
			50372: outdata = 32'd15164;
			50373: outdata = 32'd15163;
			50374: outdata = 32'd15162;
			50375: outdata = 32'd15161;
			50376: outdata = 32'd15160;
			50377: outdata = 32'd15159;
			50378: outdata = 32'd15158;
			50379: outdata = 32'd15157;
			50380: outdata = 32'd15156;
			50381: outdata = 32'd15155;
			50382: outdata = 32'd15154;
			50383: outdata = 32'd15153;
			50384: outdata = 32'd15152;
			50385: outdata = 32'd15151;
			50386: outdata = 32'd15150;
			50387: outdata = 32'd15149;
			50388: outdata = 32'd15148;
			50389: outdata = 32'd15147;
			50390: outdata = 32'd15146;
			50391: outdata = 32'd15145;
			50392: outdata = 32'd15144;
			50393: outdata = 32'd15143;
			50394: outdata = 32'd15142;
			50395: outdata = 32'd15141;
			50396: outdata = 32'd15140;
			50397: outdata = 32'd15139;
			50398: outdata = 32'd15138;
			50399: outdata = 32'd15137;
			50400: outdata = 32'd15136;
			50401: outdata = 32'd15135;
			50402: outdata = 32'd15134;
			50403: outdata = 32'd15133;
			50404: outdata = 32'd15132;
			50405: outdata = 32'd15131;
			50406: outdata = 32'd15130;
			50407: outdata = 32'd15129;
			50408: outdata = 32'd15128;
			50409: outdata = 32'd15127;
			50410: outdata = 32'd15126;
			50411: outdata = 32'd15125;
			50412: outdata = 32'd15124;
			50413: outdata = 32'd15123;
			50414: outdata = 32'd15122;
			50415: outdata = 32'd15121;
			50416: outdata = 32'd15120;
			50417: outdata = 32'd15119;
			50418: outdata = 32'd15118;
			50419: outdata = 32'd15117;
			50420: outdata = 32'd15116;
			50421: outdata = 32'd15115;
			50422: outdata = 32'd15114;
			50423: outdata = 32'd15113;
			50424: outdata = 32'd15112;
			50425: outdata = 32'd15111;
			50426: outdata = 32'd15110;
			50427: outdata = 32'd15109;
			50428: outdata = 32'd15108;
			50429: outdata = 32'd15107;
			50430: outdata = 32'd15106;
			50431: outdata = 32'd15105;
			50432: outdata = 32'd15104;
			50433: outdata = 32'd15103;
			50434: outdata = 32'd15102;
			50435: outdata = 32'd15101;
			50436: outdata = 32'd15100;
			50437: outdata = 32'd15099;
			50438: outdata = 32'd15098;
			50439: outdata = 32'd15097;
			50440: outdata = 32'd15096;
			50441: outdata = 32'd15095;
			50442: outdata = 32'd15094;
			50443: outdata = 32'd15093;
			50444: outdata = 32'd15092;
			50445: outdata = 32'd15091;
			50446: outdata = 32'd15090;
			50447: outdata = 32'd15089;
			50448: outdata = 32'd15088;
			50449: outdata = 32'd15087;
			50450: outdata = 32'd15086;
			50451: outdata = 32'd15085;
			50452: outdata = 32'd15084;
			50453: outdata = 32'd15083;
			50454: outdata = 32'd15082;
			50455: outdata = 32'd15081;
			50456: outdata = 32'd15080;
			50457: outdata = 32'd15079;
			50458: outdata = 32'd15078;
			50459: outdata = 32'd15077;
			50460: outdata = 32'd15076;
			50461: outdata = 32'd15075;
			50462: outdata = 32'd15074;
			50463: outdata = 32'd15073;
			50464: outdata = 32'd15072;
			50465: outdata = 32'd15071;
			50466: outdata = 32'd15070;
			50467: outdata = 32'd15069;
			50468: outdata = 32'd15068;
			50469: outdata = 32'd15067;
			50470: outdata = 32'd15066;
			50471: outdata = 32'd15065;
			50472: outdata = 32'd15064;
			50473: outdata = 32'd15063;
			50474: outdata = 32'd15062;
			50475: outdata = 32'd15061;
			50476: outdata = 32'd15060;
			50477: outdata = 32'd15059;
			50478: outdata = 32'd15058;
			50479: outdata = 32'd15057;
			50480: outdata = 32'd15056;
			50481: outdata = 32'd15055;
			50482: outdata = 32'd15054;
			50483: outdata = 32'd15053;
			50484: outdata = 32'd15052;
			50485: outdata = 32'd15051;
			50486: outdata = 32'd15050;
			50487: outdata = 32'd15049;
			50488: outdata = 32'd15048;
			50489: outdata = 32'd15047;
			50490: outdata = 32'd15046;
			50491: outdata = 32'd15045;
			50492: outdata = 32'd15044;
			50493: outdata = 32'd15043;
			50494: outdata = 32'd15042;
			50495: outdata = 32'd15041;
			50496: outdata = 32'd15040;
			50497: outdata = 32'd15039;
			50498: outdata = 32'd15038;
			50499: outdata = 32'd15037;
			50500: outdata = 32'd15036;
			50501: outdata = 32'd15035;
			50502: outdata = 32'd15034;
			50503: outdata = 32'd15033;
			50504: outdata = 32'd15032;
			50505: outdata = 32'd15031;
			50506: outdata = 32'd15030;
			50507: outdata = 32'd15029;
			50508: outdata = 32'd15028;
			50509: outdata = 32'd15027;
			50510: outdata = 32'd15026;
			50511: outdata = 32'd15025;
			50512: outdata = 32'd15024;
			50513: outdata = 32'd15023;
			50514: outdata = 32'd15022;
			50515: outdata = 32'd15021;
			50516: outdata = 32'd15020;
			50517: outdata = 32'd15019;
			50518: outdata = 32'd15018;
			50519: outdata = 32'd15017;
			50520: outdata = 32'd15016;
			50521: outdata = 32'd15015;
			50522: outdata = 32'd15014;
			50523: outdata = 32'd15013;
			50524: outdata = 32'd15012;
			50525: outdata = 32'd15011;
			50526: outdata = 32'd15010;
			50527: outdata = 32'd15009;
			50528: outdata = 32'd15008;
			50529: outdata = 32'd15007;
			50530: outdata = 32'd15006;
			50531: outdata = 32'd15005;
			50532: outdata = 32'd15004;
			50533: outdata = 32'd15003;
			50534: outdata = 32'd15002;
			50535: outdata = 32'd15001;
			50536: outdata = 32'd15000;
			50537: outdata = 32'd14999;
			50538: outdata = 32'd14998;
			50539: outdata = 32'd14997;
			50540: outdata = 32'd14996;
			50541: outdata = 32'd14995;
			50542: outdata = 32'd14994;
			50543: outdata = 32'd14993;
			50544: outdata = 32'd14992;
			50545: outdata = 32'd14991;
			50546: outdata = 32'd14990;
			50547: outdata = 32'd14989;
			50548: outdata = 32'd14988;
			50549: outdata = 32'd14987;
			50550: outdata = 32'd14986;
			50551: outdata = 32'd14985;
			50552: outdata = 32'd14984;
			50553: outdata = 32'd14983;
			50554: outdata = 32'd14982;
			50555: outdata = 32'd14981;
			50556: outdata = 32'd14980;
			50557: outdata = 32'd14979;
			50558: outdata = 32'd14978;
			50559: outdata = 32'd14977;
			50560: outdata = 32'd14976;
			50561: outdata = 32'd14975;
			50562: outdata = 32'd14974;
			50563: outdata = 32'd14973;
			50564: outdata = 32'd14972;
			50565: outdata = 32'd14971;
			50566: outdata = 32'd14970;
			50567: outdata = 32'd14969;
			50568: outdata = 32'd14968;
			50569: outdata = 32'd14967;
			50570: outdata = 32'd14966;
			50571: outdata = 32'd14965;
			50572: outdata = 32'd14964;
			50573: outdata = 32'd14963;
			50574: outdata = 32'd14962;
			50575: outdata = 32'd14961;
			50576: outdata = 32'd14960;
			50577: outdata = 32'd14959;
			50578: outdata = 32'd14958;
			50579: outdata = 32'd14957;
			50580: outdata = 32'd14956;
			50581: outdata = 32'd14955;
			50582: outdata = 32'd14954;
			50583: outdata = 32'd14953;
			50584: outdata = 32'd14952;
			50585: outdata = 32'd14951;
			50586: outdata = 32'd14950;
			50587: outdata = 32'd14949;
			50588: outdata = 32'd14948;
			50589: outdata = 32'd14947;
			50590: outdata = 32'd14946;
			50591: outdata = 32'd14945;
			50592: outdata = 32'd14944;
			50593: outdata = 32'd14943;
			50594: outdata = 32'd14942;
			50595: outdata = 32'd14941;
			50596: outdata = 32'd14940;
			50597: outdata = 32'd14939;
			50598: outdata = 32'd14938;
			50599: outdata = 32'd14937;
			50600: outdata = 32'd14936;
			50601: outdata = 32'd14935;
			50602: outdata = 32'd14934;
			50603: outdata = 32'd14933;
			50604: outdata = 32'd14932;
			50605: outdata = 32'd14931;
			50606: outdata = 32'd14930;
			50607: outdata = 32'd14929;
			50608: outdata = 32'd14928;
			50609: outdata = 32'd14927;
			50610: outdata = 32'd14926;
			50611: outdata = 32'd14925;
			50612: outdata = 32'd14924;
			50613: outdata = 32'd14923;
			50614: outdata = 32'd14922;
			50615: outdata = 32'd14921;
			50616: outdata = 32'd14920;
			50617: outdata = 32'd14919;
			50618: outdata = 32'd14918;
			50619: outdata = 32'd14917;
			50620: outdata = 32'd14916;
			50621: outdata = 32'd14915;
			50622: outdata = 32'd14914;
			50623: outdata = 32'd14913;
			50624: outdata = 32'd14912;
			50625: outdata = 32'd14911;
			50626: outdata = 32'd14910;
			50627: outdata = 32'd14909;
			50628: outdata = 32'd14908;
			50629: outdata = 32'd14907;
			50630: outdata = 32'd14906;
			50631: outdata = 32'd14905;
			50632: outdata = 32'd14904;
			50633: outdata = 32'd14903;
			50634: outdata = 32'd14902;
			50635: outdata = 32'd14901;
			50636: outdata = 32'd14900;
			50637: outdata = 32'd14899;
			50638: outdata = 32'd14898;
			50639: outdata = 32'd14897;
			50640: outdata = 32'd14896;
			50641: outdata = 32'd14895;
			50642: outdata = 32'd14894;
			50643: outdata = 32'd14893;
			50644: outdata = 32'd14892;
			50645: outdata = 32'd14891;
			50646: outdata = 32'd14890;
			50647: outdata = 32'd14889;
			50648: outdata = 32'd14888;
			50649: outdata = 32'd14887;
			50650: outdata = 32'd14886;
			50651: outdata = 32'd14885;
			50652: outdata = 32'd14884;
			50653: outdata = 32'd14883;
			50654: outdata = 32'd14882;
			50655: outdata = 32'd14881;
			50656: outdata = 32'd14880;
			50657: outdata = 32'd14879;
			50658: outdata = 32'd14878;
			50659: outdata = 32'd14877;
			50660: outdata = 32'd14876;
			50661: outdata = 32'd14875;
			50662: outdata = 32'd14874;
			50663: outdata = 32'd14873;
			50664: outdata = 32'd14872;
			50665: outdata = 32'd14871;
			50666: outdata = 32'd14870;
			50667: outdata = 32'd14869;
			50668: outdata = 32'd14868;
			50669: outdata = 32'd14867;
			50670: outdata = 32'd14866;
			50671: outdata = 32'd14865;
			50672: outdata = 32'd14864;
			50673: outdata = 32'd14863;
			50674: outdata = 32'd14862;
			50675: outdata = 32'd14861;
			50676: outdata = 32'd14860;
			50677: outdata = 32'd14859;
			50678: outdata = 32'd14858;
			50679: outdata = 32'd14857;
			50680: outdata = 32'd14856;
			50681: outdata = 32'd14855;
			50682: outdata = 32'd14854;
			50683: outdata = 32'd14853;
			50684: outdata = 32'd14852;
			50685: outdata = 32'd14851;
			50686: outdata = 32'd14850;
			50687: outdata = 32'd14849;
			50688: outdata = 32'd14848;
			50689: outdata = 32'd14847;
			50690: outdata = 32'd14846;
			50691: outdata = 32'd14845;
			50692: outdata = 32'd14844;
			50693: outdata = 32'd14843;
			50694: outdata = 32'd14842;
			50695: outdata = 32'd14841;
			50696: outdata = 32'd14840;
			50697: outdata = 32'd14839;
			50698: outdata = 32'd14838;
			50699: outdata = 32'd14837;
			50700: outdata = 32'd14836;
			50701: outdata = 32'd14835;
			50702: outdata = 32'd14834;
			50703: outdata = 32'd14833;
			50704: outdata = 32'd14832;
			50705: outdata = 32'd14831;
			50706: outdata = 32'd14830;
			50707: outdata = 32'd14829;
			50708: outdata = 32'd14828;
			50709: outdata = 32'd14827;
			50710: outdata = 32'd14826;
			50711: outdata = 32'd14825;
			50712: outdata = 32'd14824;
			50713: outdata = 32'd14823;
			50714: outdata = 32'd14822;
			50715: outdata = 32'd14821;
			50716: outdata = 32'd14820;
			50717: outdata = 32'd14819;
			50718: outdata = 32'd14818;
			50719: outdata = 32'd14817;
			50720: outdata = 32'd14816;
			50721: outdata = 32'd14815;
			50722: outdata = 32'd14814;
			50723: outdata = 32'd14813;
			50724: outdata = 32'd14812;
			50725: outdata = 32'd14811;
			50726: outdata = 32'd14810;
			50727: outdata = 32'd14809;
			50728: outdata = 32'd14808;
			50729: outdata = 32'd14807;
			50730: outdata = 32'd14806;
			50731: outdata = 32'd14805;
			50732: outdata = 32'd14804;
			50733: outdata = 32'd14803;
			50734: outdata = 32'd14802;
			50735: outdata = 32'd14801;
			50736: outdata = 32'd14800;
			50737: outdata = 32'd14799;
			50738: outdata = 32'd14798;
			50739: outdata = 32'd14797;
			50740: outdata = 32'd14796;
			50741: outdata = 32'd14795;
			50742: outdata = 32'd14794;
			50743: outdata = 32'd14793;
			50744: outdata = 32'd14792;
			50745: outdata = 32'd14791;
			50746: outdata = 32'd14790;
			50747: outdata = 32'd14789;
			50748: outdata = 32'd14788;
			50749: outdata = 32'd14787;
			50750: outdata = 32'd14786;
			50751: outdata = 32'd14785;
			50752: outdata = 32'd14784;
			50753: outdata = 32'd14783;
			50754: outdata = 32'd14782;
			50755: outdata = 32'd14781;
			50756: outdata = 32'd14780;
			50757: outdata = 32'd14779;
			50758: outdata = 32'd14778;
			50759: outdata = 32'd14777;
			50760: outdata = 32'd14776;
			50761: outdata = 32'd14775;
			50762: outdata = 32'd14774;
			50763: outdata = 32'd14773;
			50764: outdata = 32'd14772;
			50765: outdata = 32'd14771;
			50766: outdata = 32'd14770;
			50767: outdata = 32'd14769;
			50768: outdata = 32'd14768;
			50769: outdata = 32'd14767;
			50770: outdata = 32'd14766;
			50771: outdata = 32'd14765;
			50772: outdata = 32'd14764;
			50773: outdata = 32'd14763;
			50774: outdata = 32'd14762;
			50775: outdata = 32'd14761;
			50776: outdata = 32'd14760;
			50777: outdata = 32'd14759;
			50778: outdata = 32'd14758;
			50779: outdata = 32'd14757;
			50780: outdata = 32'd14756;
			50781: outdata = 32'd14755;
			50782: outdata = 32'd14754;
			50783: outdata = 32'd14753;
			50784: outdata = 32'd14752;
			50785: outdata = 32'd14751;
			50786: outdata = 32'd14750;
			50787: outdata = 32'd14749;
			50788: outdata = 32'd14748;
			50789: outdata = 32'd14747;
			50790: outdata = 32'd14746;
			50791: outdata = 32'd14745;
			50792: outdata = 32'd14744;
			50793: outdata = 32'd14743;
			50794: outdata = 32'd14742;
			50795: outdata = 32'd14741;
			50796: outdata = 32'd14740;
			50797: outdata = 32'd14739;
			50798: outdata = 32'd14738;
			50799: outdata = 32'd14737;
			50800: outdata = 32'd14736;
			50801: outdata = 32'd14735;
			50802: outdata = 32'd14734;
			50803: outdata = 32'd14733;
			50804: outdata = 32'd14732;
			50805: outdata = 32'd14731;
			50806: outdata = 32'd14730;
			50807: outdata = 32'd14729;
			50808: outdata = 32'd14728;
			50809: outdata = 32'd14727;
			50810: outdata = 32'd14726;
			50811: outdata = 32'd14725;
			50812: outdata = 32'd14724;
			50813: outdata = 32'd14723;
			50814: outdata = 32'd14722;
			50815: outdata = 32'd14721;
			50816: outdata = 32'd14720;
			50817: outdata = 32'd14719;
			50818: outdata = 32'd14718;
			50819: outdata = 32'd14717;
			50820: outdata = 32'd14716;
			50821: outdata = 32'd14715;
			50822: outdata = 32'd14714;
			50823: outdata = 32'd14713;
			50824: outdata = 32'd14712;
			50825: outdata = 32'd14711;
			50826: outdata = 32'd14710;
			50827: outdata = 32'd14709;
			50828: outdata = 32'd14708;
			50829: outdata = 32'd14707;
			50830: outdata = 32'd14706;
			50831: outdata = 32'd14705;
			50832: outdata = 32'd14704;
			50833: outdata = 32'd14703;
			50834: outdata = 32'd14702;
			50835: outdata = 32'd14701;
			50836: outdata = 32'd14700;
			50837: outdata = 32'd14699;
			50838: outdata = 32'd14698;
			50839: outdata = 32'd14697;
			50840: outdata = 32'd14696;
			50841: outdata = 32'd14695;
			50842: outdata = 32'd14694;
			50843: outdata = 32'd14693;
			50844: outdata = 32'd14692;
			50845: outdata = 32'd14691;
			50846: outdata = 32'd14690;
			50847: outdata = 32'd14689;
			50848: outdata = 32'd14688;
			50849: outdata = 32'd14687;
			50850: outdata = 32'd14686;
			50851: outdata = 32'd14685;
			50852: outdata = 32'd14684;
			50853: outdata = 32'd14683;
			50854: outdata = 32'd14682;
			50855: outdata = 32'd14681;
			50856: outdata = 32'd14680;
			50857: outdata = 32'd14679;
			50858: outdata = 32'd14678;
			50859: outdata = 32'd14677;
			50860: outdata = 32'd14676;
			50861: outdata = 32'd14675;
			50862: outdata = 32'd14674;
			50863: outdata = 32'd14673;
			50864: outdata = 32'd14672;
			50865: outdata = 32'd14671;
			50866: outdata = 32'd14670;
			50867: outdata = 32'd14669;
			50868: outdata = 32'd14668;
			50869: outdata = 32'd14667;
			50870: outdata = 32'd14666;
			50871: outdata = 32'd14665;
			50872: outdata = 32'd14664;
			50873: outdata = 32'd14663;
			50874: outdata = 32'd14662;
			50875: outdata = 32'd14661;
			50876: outdata = 32'd14660;
			50877: outdata = 32'd14659;
			50878: outdata = 32'd14658;
			50879: outdata = 32'd14657;
			50880: outdata = 32'd14656;
			50881: outdata = 32'd14655;
			50882: outdata = 32'd14654;
			50883: outdata = 32'd14653;
			50884: outdata = 32'd14652;
			50885: outdata = 32'd14651;
			50886: outdata = 32'd14650;
			50887: outdata = 32'd14649;
			50888: outdata = 32'd14648;
			50889: outdata = 32'd14647;
			50890: outdata = 32'd14646;
			50891: outdata = 32'd14645;
			50892: outdata = 32'd14644;
			50893: outdata = 32'd14643;
			50894: outdata = 32'd14642;
			50895: outdata = 32'd14641;
			50896: outdata = 32'd14640;
			50897: outdata = 32'd14639;
			50898: outdata = 32'd14638;
			50899: outdata = 32'd14637;
			50900: outdata = 32'd14636;
			50901: outdata = 32'd14635;
			50902: outdata = 32'd14634;
			50903: outdata = 32'd14633;
			50904: outdata = 32'd14632;
			50905: outdata = 32'd14631;
			50906: outdata = 32'd14630;
			50907: outdata = 32'd14629;
			50908: outdata = 32'd14628;
			50909: outdata = 32'd14627;
			50910: outdata = 32'd14626;
			50911: outdata = 32'd14625;
			50912: outdata = 32'd14624;
			50913: outdata = 32'd14623;
			50914: outdata = 32'd14622;
			50915: outdata = 32'd14621;
			50916: outdata = 32'd14620;
			50917: outdata = 32'd14619;
			50918: outdata = 32'd14618;
			50919: outdata = 32'd14617;
			50920: outdata = 32'd14616;
			50921: outdata = 32'd14615;
			50922: outdata = 32'd14614;
			50923: outdata = 32'd14613;
			50924: outdata = 32'd14612;
			50925: outdata = 32'd14611;
			50926: outdata = 32'd14610;
			50927: outdata = 32'd14609;
			50928: outdata = 32'd14608;
			50929: outdata = 32'd14607;
			50930: outdata = 32'd14606;
			50931: outdata = 32'd14605;
			50932: outdata = 32'd14604;
			50933: outdata = 32'd14603;
			50934: outdata = 32'd14602;
			50935: outdata = 32'd14601;
			50936: outdata = 32'd14600;
			50937: outdata = 32'd14599;
			50938: outdata = 32'd14598;
			50939: outdata = 32'd14597;
			50940: outdata = 32'd14596;
			50941: outdata = 32'd14595;
			50942: outdata = 32'd14594;
			50943: outdata = 32'd14593;
			50944: outdata = 32'd14592;
			50945: outdata = 32'd14591;
			50946: outdata = 32'd14590;
			50947: outdata = 32'd14589;
			50948: outdata = 32'd14588;
			50949: outdata = 32'd14587;
			50950: outdata = 32'd14586;
			50951: outdata = 32'd14585;
			50952: outdata = 32'd14584;
			50953: outdata = 32'd14583;
			50954: outdata = 32'd14582;
			50955: outdata = 32'd14581;
			50956: outdata = 32'd14580;
			50957: outdata = 32'd14579;
			50958: outdata = 32'd14578;
			50959: outdata = 32'd14577;
			50960: outdata = 32'd14576;
			50961: outdata = 32'd14575;
			50962: outdata = 32'd14574;
			50963: outdata = 32'd14573;
			50964: outdata = 32'd14572;
			50965: outdata = 32'd14571;
			50966: outdata = 32'd14570;
			50967: outdata = 32'd14569;
			50968: outdata = 32'd14568;
			50969: outdata = 32'd14567;
			50970: outdata = 32'd14566;
			50971: outdata = 32'd14565;
			50972: outdata = 32'd14564;
			50973: outdata = 32'd14563;
			50974: outdata = 32'd14562;
			50975: outdata = 32'd14561;
			50976: outdata = 32'd14560;
			50977: outdata = 32'd14559;
			50978: outdata = 32'd14558;
			50979: outdata = 32'd14557;
			50980: outdata = 32'd14556;
			50981: outdata = 32'd14555;
			50982: outdata = 32'd14554;
			50983: outdata = 32'd14553;
			50984: outdata = 32'd14552;
			50985: outdata = 32'd14551;
			50986: outdata = 32'd14550;
			50987: outdata = 32'd14549;
			50988: outdata = 32'd14548;
			50989: outdata = 32'd14547;
			50990: outdata = 32'd14546;
			50991: outdata = 32'd14545;
			50992: outdata = 32'd14544;
			50993: outdata = 32'd14543;
			50994: outdata = 32'd14542;
			50995: outdata = 32'd14541;
			50996: outdata = 32'd14540;
			50997: outdata = 32'd14539;
			50998: outdata = 32'd14538;
			50999: outdata = 32'd14537;
			51000: outdata = 32'd14536;
			51001: outdata = 32'd14535;
			51002: outdata = 32'd14534;
			51003: outdata = 32'd14533;
			51004: outdata = 32'd14532;
			51005: outdata = 32'd14531;
			51006: outdata = 32'd14530;
			51007: outdata = 32'd14529;
			51008: outdata = 32'd14528;
			51009: outdata = 32'd14527;
			51010: outdata = 32'd14526;
			51011: outdata = 32'd14525;
			51012: outdata = 32'd14524;
			51013: outdata = 32'd14523;
			51014: outdata = 32'd14522;
			51015: outdata = 32'd14521;
			51016: outdata = 32'd14520;
			51017: outdata = 32'd14519;
			51018: outdata = 32'd14518;
			51019: outdata = 32'd14517;
			51020: outdata = 32'd14516;
			51021: outdata = 32'd14515;
			51022: outdata = 32'd14514;
			51023: outdata = 32'd14513;
			51024: outdata = 32'd14512;
			51025: outdata = 32'd14511;
			51026: outdata = 32'd14510;
			51027: outdata = 32'd14509;
			51028: outdata = 32'd14508;
			51029: outdata = 32'd14507;
			51030: outdata = 32'd14506;
			51031: outdata = 32'd14505;
			51032: outdata = 32'd14504;
			51033: outdata = 32'd14503;
			51034: outdata = 32'd14502;
			51035: outdata = 32'd14501;
			51036: outdata = 32'd14500;
			51037: outdata = 32'd14499;
			51038: outdata = 32'd14498;
			51039: outdata = 32'd14497;
			51040: outdata = 32'd14496;
			51041: outdata = 32'd14495;
			51042: outdata = 32'd14494;
			51043: outdata = 32'd14493;
			51044: outdata = 32'd14492;
			51045: outdata = 32'd14491;
			51046: outdata = 32'd14490;
			51047: outdata = 32'd14489;
			51048: outdata = 32'd14488;
			51049: outdata = 32'd14487;
			51050: outdata = 32'd14486;
			51051: outdata = 32'd14485;
			51052: outdata = 32'd14484;
			51053: outdata = 32'd14483;
			51054: outdata = 32'd14482;
			51055: outdata = 32'd14481;
			51056: outdata = 32'd14480;
			51057: outdata = 32'd14479;
			51058: outdata = 32'd14478;
			51059: outdata = 32'd14477;
			51060: outdata = 32'd14476;
			51061: outdata = 32'd14475;
			51062: outdata = 32'd14474;
			51063: outdata = 32'd14473;
			51064: outdata = 32'd14472;
			51065: outdata = 32'd14471;
			51066: outdata = 32'd14470;
			51067: outdata = 32'd14469;
			51068: outdata = 32'd14468;
			51069: outdata = 32'd14467;
			51070: outdata = 32'd14466;
			51071: outdata = 32'd14465;
			51072: outdata = 32'd14464;
			51073: outdata = 32'd14463;
			51074: outdata = 32'd14462;
			51075: outdata = 32'd14461;
			51076: outdata = 32'd14460;
			51077: outdata = 32'd14459;
			51078: outdata = 32'd14458;
			51079: outdata = 32'd14457;
			51080: outdata = 32'd14456;
			51081: outdata = 32'd14455;
			51082: outdata = 32'd14454;
			51083: outdata = 32'd14453;
			51084: outdata = 32'd14452;
			51085: outdata = 32'd14451;
			51086: outdata = 32'd14450;
			51087: outdata = 32'd14449;
			51088: outdata = 32'd14448;
			51089: outdata = 32'd14447;
			51090: outdata = 32'd14446;
			51091: outdata = 32'd14445;
			51092: outdata = 32'd14444;
			51093: outdata = 32'd14443;
			51094: outdata = 32'd14442;
			51095: outdata = 32'd14441;
			51096: outdata = 32'd14440;
			51097: outdata = 32'd14439;
			51098: outdata = 32'd14438;
			51099: outdata = 32'd14437;
			51100: outdata = 32'd14436;
			51101: outdata = 32'd14435;
			51102: outdata = 32'd14434;
			51103: outdata = 32'd14433;
			51104: outdata = 32'd14432;
			51105: outdata = 32'd14431;
			51106: outdata = 32'd14430;
			51107: outdata = 32'd14429;
			51108: outdata = 32'd14428;
			51109: outdata = 32'd14427;
			51110: outdata = 32'd14426;
			51111: outdata = 32'd14425;
			51112: outdata = 32'd14424;
			51113: outdata = 32'd14423;
			51114: outdata = 32'd14422;
			51115: outdata = 32'd14421;
			51116: outdata = 32'd14420;
			51117: outdata = 32'd14419;
			51118: outdata = 32'd14418;
			51119: outdata = 32'd14417;
			51120: outdata = 32'd14416;
			51121: outdata = 32'd14415;
			51122: outdata = 32'd14414;
			51123: outdata = 32'd14413;
			51124: outdata = 32'd14412;
			51125: outdata = 32'd14411;
			51126: outdata = 32'd14410;
			51127: outdata = 32'd14409;
			51128: outdata = 32'd14408;
			51129: outdata = 32'd14407;
			51130: outdata = 32'd14406;
			51131: outdata = 32'd14405;
			51132: outdata = 32'd14404;
			51133: outdata = 32'd14403;
			51134: outdata = 32'd14402;
			51135: outdata = 32'd14401;
			51136: outdata = 32'd14400;
			51137: outdata = 32'd14399;
			51138: outdata = 32'd14398;
			51139: outdata = 32'd14397;
			51140: outdata = 32'd14396;
			51141: outdata = 32'd14395;
			51142: outdata = 32'd14394;
			51143: outdata = 32'd14393;
			51144: outdata = 32'd14392;
			51145: outdata = 32'd14391;
			51146: outdata = 32'd14390;
			51147: outdata = 32'd14389;
			51148: outdata = 32'd14388;
			51149: outdata = 32'd14387;
			51150: outdata = 32'd14386;
			51151: outdata = 32'd14385;
			51152: outdata = 32'd14384;
			51153: outdata = 32'd14383;
			51154: outdata = 32'd14382;
			51155: outdata = 32'd14381;
			51156: outdata = 32'd14380;
			51157: outdata = 32'd14379;
			51158: outdata = 32'd14378;
			51159: outdata = 32'd14377;
			51160: outdata = 32'd14376;
			51161: outdata = 32'd14375;
			51162: outdata = 32'd14374;
			51163: outdata = 32'd14373;
			51164: outdata = 32'd14372;
			51165: outdata = 32'd14371;
			51166: outdata = 32'd14370;
			51167: outdata = 32'd14369;
			51168: outdata = 32'd14368;
			51169: outdata = 32'd14367;
			51170: outdata = 32'd14366;
			51171: outdata = 32'd14365;
			51172: outdata = 32'd14364;
			51173: outdata = 32'd14363;
			51174: outdata = 32'd14362;
			51175: outdata = 32'd14361;
			51176: outdata = 32'd14360;
			51177: outdata = 32'd14359;
			51178: outdata = 32'd14358;
			51179: outdata = 32'd14357;
			51180: outdata = 32'd14356;
			51181: outdata = 32'd14355;
			51182: outdata = 32'd14354;
			51183: outdata = 32'd14353;
			51184: outdata = 32'd14352;
			51185: outdata = 32'd14351;
			51186: outdata = 32'd14350;
			51187: outdata = 32'd14349;
			51188: outdata = 32'd14348;
			51189: outdata = 32'd14347;
			51190: outdata = 32'd14346;
			51191: outdata = 32'd14345;
			51192: outdata = 32'd14344;
			51193: outdata = 32'd14343;
			51194: outdata = 32'd14342;
			51195: outdata = 32'd14341;
			51196: outdata = 32'd14340;
			51197: outdata = 32'd14339;
			51198: outdata = 32'd14338;
			51199: outdata = 32'd14337;
			51200: outdata = 32'd14336;
			51201: outdata = 32'd14335;
			51202: outdata = 32'd14334;
			51203: outdata = 32'd14333;
			51204: outdata = 32'd14332;
			51205: outdata = 32'd14331;
			51206: outdata = 32'd14330;
			51207: outdata = 32'd14329;
			51208: outdata = 32'd14328;
			51209: outdata = 32'd14327;
			51210: outdata = 32'd14326;
			51211: outdata = 32'd14325;
			51212: outdata = 32'd14324;
			51213: outdata = 32'd14323;
			51214: outdata = 32'd14322;
			51215: outdata = 32'd14321;
			51216: outdata = 32'd14320;
			51217: outdata = 32'd14319;
			51218: outdata = 32'd14318;
			51219: outdata = 32'd14317;
			51220: outdata = 32'd14316;
			51221: outdata = 32'd14315;
			51222: outdata = 32'd14314;
			51223: outdata = 32'd14313;
			51224: outdata = 32'd14312;
			51225: outdata = 32'd14311;
			51226: outdata = 32'd14310;
			51227: outdata = 32'd14309;
			51228: outdata = 32'd14308;
			51229: outdata = 32'd14307;
			51230: outdata = 32'd14306;
			51231: outdata = 32'd14305;
			51232: outdata = 32'd14304;
			51233: outdata = 32'd14303;
			51234: outdata = 32'd14302;
			51235: outdata = 32'd14301;
			51236: outdata = 32'd14300;
			51237: outdata = 32'd14299;
			51238: outdata = 32'd14298;
			51239: outdata = 32'd14297;
			51240: outdata = 32'd14296;
			51241: outdata = 32'd14295;
			51242: outdata = 32'd14294;
			51243: outdata = 32'd14293;
			51244: outdata = 32'd14292;
			51245: outdata = 32'd14291;
			51246: outdata = 32'd14290;
			51247: outdata = 32'd14289;
			51248: outdata = 32'd14288;
			51249: outdata = 32'd14287;
			51250: outdata = 32'd14286;
			51251: outdata = 32'd14285;
			51252: outdata = 32'd14284;
			51253: outdata = 32'd14283;
			51254: outdata = 32'd14282;
			51255: outdata = 32'd14281;
			51256: outdata = 32'd14280;
			51257: outdata = 32'd14279;
			51258: outdata = 32'd14278;
			51259: outdata = 32'd14277;
			51260: outdata = 32'd14276;
			51261: outdata = 32'd14275;
			51262: outdata = 32'd14274;
			51263: outdata = 32'd14273;
			51264: outdata = 32'd14272;
			51265: outdata = 32'd14271;
			51266: outdata = 32'd14270;
			51267: outdata = 32'd14269;
			51268: outdata = 32'd14268;
			51269: outdata = 32'd14267;
			51270: outdata = 32'd14266;
			51271: outdata = 32'd14265;
			51272: outdata = 32'd14264;
			51273: outdata = 32'd14263;
			51274: outdata = 32'd14262;
			51275: outdata = 32'd14261;
			51276: outdata = 32'd14260;
			51277: outdata = 32'd14259;
			51278: outdata = 32'd14258;
			51279: outdata = 32'd14257;
			51280: outdata = 32'd14256;
			51281: outdata = 32'd14255;
			51282: outdata = 32'd14254;
			51283: outdata = 32'd14253;
			51284: outdata = 32'd14252;
			51285: outdata = 32'd14251;
			51286: outdata = 32'd14250;
			51287: outdata = 32'd14249;
			51288: outdata = 32'd14248;
			51289: outdata = 32'd14247;
			51290: outdata = 32'd14246;
			51291: outdata = 32'd14245;
			51292: outdata = 32'd14244;
			51293: outdata = 32'd14243;
			51294: outdata = 32'd14242;
			51295: outdata = 32'd14241;
			51296: outdata = 32'd14240;
			51297: outdata = 32'd14239;
			51298: outdata = 32'd14238;
			51299: outdata = 32'd14237;
			51300: outdata = 32'd14236;
			51301: outdata = 32'd14235;
			51302: outdata = 32'd14234;
			51303: outdata = 32'd14233;
			51304: outdata = 32'd14232;
			51305: outdata = 32'd14231;
			51306: outdata = 32'd14230;
			51307: outdata = 32'd14229;
			51308: outdata = 32'd14228;
			51309: outdata = 32'd14227;
			51310: outdata = 32'd14226;
			51311: outdata = 32'd14225;
			51312: outdata = 32'd14224;
			51313: outdata = 32'd14223;
			51314: outdata = 32'd14222;
			51315: outdata = 32'd14221;
			51316: outdata = 32'd14220;
			51317: outdata = 32'd14219;
			51318: outdata = 32'd14218;
			51319: outdata = 32'd14217;
			51320: outdata = 32'd14216;
			51321: outdata = 32'd14215;
			51322: outdata = 32'd14214;
			51323: outdata = 32'd14213;
			51324: outdata = 32'd14212;
			51325: outdata = 32'd14211;
			51326: outdata = 32'd14210;
			51327: outdata = 32'd14209;
			51328: outdata = 32'd14208;
			51329: outdata = 32'd14207;
			51330: outdata = 32'd14206;
			51331: outdata = 32'd14205;
			51332: outdata = 32'd14204;
			51333: outdata = 32'd14203;
			51334: outdata = 32'd14202;
			51335: outdata = 32'd14201;
			51336: outdata = 32'd14200;
			51337: outdata = 32'd14199;
			51338: outdata = 32'd14198;
			51339: outdata = 32'd14197;
			51340: outdata = 32'd14196;
			51341: outdata = 32'd14195;
			51342: outdata = 32'd14194;
			51343: outdata = 32'd14193;
			51344: outdata = 32'd14192;
			51345: outdata = 32'd14191;
			51346: outdata = 32'd14190;
			51347: outdata = 32'd14189;
			51348: outdata = 32'd14188;
			51349: outdata = 32'd14187;
			51350: outdata = 32'd14186;
			51351: outdata = 32'd14185;
			51352: outdata = 32'd14184;
			51353: outdata = 32'd14183;
			51354: outdata = 32'd14182;
			51355: outdata = 32'd14181;
			51356: outdata = 32'd14180;
			51357: outdata = 32'd14179;
			51358: outdata = 32'd14178;
			51359: outdata = 32'd14177;
			51360: outdata = 32'd14176;
			51361: outdata = 32'd14175;
			51362: outdata = 32'd14174;
			51363: outdata = 32'd14173;
			51364: outdata = 32'd14172;
			51365: outdata = 32'd14171;
			51366: outdata = 32'd14170;
			51367: outdata = 32'd14169;
			51368: outdata = 32'd14168;
			51369: outdata = 32'd14167;
			51370: outdata = 32'd14166;
			51371: outdata = 32'd14165;
			51372: outdata = 32'd14164;
			51373: outdata = 32'd14163;
			51374: outdata = 32'd14162;
			51375: outdata = 32'd14161;
			51376: outdata = 32'd14160;
			51377: outdata = 32'd14159;
			51378: outdata = 32'd14158;
			51379: outdata = 32'd14157;
			51380: outdata = 32'd14156;
			51381: outdata = 32'd14155;
			51382: outdata = 32'd14154;
			51383: outdata = 32'd14153;
			51384: outdata = 32'd14152;
			51385: outdata = 32'd14151;
			51386: outdata = 32'd14150;
			51387: outdata = 32'd14149;
			51388: outdata = 32'd14148;
			51389: outdata = 32'd14147;
			51390: outdata = 32'd14146;
			51391: outdata = 32'd14145;
			51392: outdata = 32'd14144;
			51393: outdata = 32'd14143;
			51394: outdata = 32'd14142;
			51395: outdata = 32'd14141;
			51396: outdata = 32'd14140;
			51397: outdata = 32'd14139;
			51398: outdata = 32'd14138;
			51399: outdata = 32'd14137;
			51400: outdata = 32'd14136;
			51401: outdata = 32'd14135;
			51402: outdata = 32'd14134;
			51403: outdata = 32'd14133;
			51404: outdata = 32'd14132;
			51405: outdata = 32'd14131;
			51406: outdata = 32'd14130;
			51407: outdata = 32'd14129;
			51408: outdata = 32'd14128;
			51409: outdata = 32'd14127;
			51410: outdata = 32'd14126;
			51411: outdata = 32'd14125;
			51412: outdata = 32'd14124;
			51413: outdata = 32'd14123;
			51414: outdata = 32'd14122;
			51415: outdata = 32'd14121;
			51416: outdata = 32'd14120;
			51417: outdata = 32'd14119;
			51418: outdata = 32'd14118;
			51419: outdata = 32'd14117;
			51420: outdata = 32'd14116;
			51421: outdata = 32'd14115;
			51422: outdata = 32'd14114;
			51423: outdata = 32'd14113;
			51424: outdata = 32'd14112;
			51425: outdata = 32'd14111;
			51426: outdata = 32'd14110;
			51427: outdata = 32'd14109;
			51428: outdata = 32'd14108;
			51429: outdata = 32'd14107;
			51430: outdata = 32'd14106;
			51431: outdata = 32'd14105;
			51432: outdata = 32'd14104;
			51433: outdata = 32'd14103;
			51434: outdata = 32'd14102;
			51435: outdata = 32'd14101;
			51436: outdata = 32'd14100;
			51437: outdata = 32'd14099;
			51438: outdata = 32'd14098;
			51439: outdata = 32'd14097;
			51440: outdata = 32'd14096;
			51441: outdata = 32'd14095;
			51442: outdata = 32'd14094;
			51443: outdata = 32'd14093;
			51444: outdata = 32'd14092;
			51445: outdata = 32'd14091;
			51446: outdata = 32'd14090;
			51447: outdata = 32'd14089;
			51448: outdata = 32'd14088;
			51449: outdata = 32'd14087;
			51450: outdata = 32'd14086;
			51451: outdata = 32'd14085;
			51452: outdata = 32'd14084;
			51453: outdata = 32'd14083;
			51454: outdata = 32'd14082;
			51455: outdata = 32'd14081;
			51456: outdata = 32'd14080;
			51457: outdata = 32'd14079;
			51458: outdata = 32'd14078;
			51459: outdata = 32'd14077;
			51460: outdata = 32'd14076;
			51461: outdata = 32'd14075;
			51462: outdata = 32'd14074;
			51463: outdata = 32'd14073;
			51464: outdata = 32'd14072;
			51465: outdata = 32'd14071;
			51466: outdata = 32'd14070;
			51467: outdata = 32'd14069;
			51468: outdata = 32'd14068;
			51469: outdata = 32'd14067;
			51470: outdata = 32'd14066;
			51471: outdata = 32'd14065;
			51472: outdata = 32'd14064;
			51473: outdata = 32'd14063;
			51474: outdata = 32'd14062;
			51475: outdata = 32'd14061;
			51476: outdata = 32'd14060;
			51477: outdata = 32'd14059;
			51478: outdata = 32'd14058;
			51479: outdata = 32'd14057;
			51480: outdata = 32'd14056;
			51481: outdata = 32'd14055;
			51482: outdata = 32'd14054;
			51483: outdata = 32'd14053;
			51484: outdata = 32'd14052;
			51485: outdata = 32'd14051;
			51486: outdata = 32'd14050;
			51487: outdata = 32'd14049;
			51488: outdata = 32'd14048;
			51489: outdata = 32'd14047;
			51490: outdata = 32'd14046;
			51491: outdata = 32'd14045;
			51492: outdata = 32'd14044;
			51493: outdata = 32'd14043;
			51494: outdata = 32'd14042;
			51495: outdata = 32'd14041;
			51496: outdata = 32'd14040;
			51497: outdata = 32'd14039;
			51498: outdata = 32'd14038;
			51499: outdata = 32'd14037;
			51500: outdata = 32'd14036;
			51501: outdata = 32'd14035;
			51502: outdata = 32'd14034;
			51503: outdata = 32'd14033;
			51504: outdata = 32'd14032;
			51505: outdata = 32'd14031;
			51506: outdata = 32'd14030;
			51507: outdata = 32'd14029;
			51508: outdata = 32'd14028;
			51509: outdata = 32'd14027;
			51510: outdata = 32'd14026;
			51511: outdata = 32'd14025;
			51512: outdata = 32'd14024;
			51513: outdata = 32'd14023;
			51514: outdata = 32'd14022;
			51515: outdata = 32'd14021;
			51516: outdata = 32'd14020;
			51517: outdata = 32'd14019;
			51518: outdata = 32'd14018;
			51519: outdata = 32'd14017;
			51520: outdata = 32'd14016;
			51521: outdata = 32'd14015;
			51522: outdata = 32'd14014;
			51523: outdata = 32'd14013;
			51524: outdata = 32'd14012;
			51525: outdata = 32'd14011;
			51526: outdata = 32'd14010;
			51527: outdata = 32'd14009;
			51528: outdata = 32'd14008;
			51529: outdata = 32'd14007;
			51530: outdata = 32'd14006;
			51531: outdata = 32'd14005;
			51532: outdata = 32'd14004;
			51533: outdata = 32'd14003;
			51534: outdata = 32'd14002;
			51535: outdata = 32'd14001;
			51536: outdata = 32'd14000;
			51537: outdata = 32'd13999;
			51538: outdata = 32'd13998;
			51539: outdata = 32'd13997;
			51540: outdata = 32'd13996;
			51541: outdata = 32'd13995;
			51542: outdata = 32'd13994;
			51543: outdata = 32'd13993;
			51544: outdata = 32'd13992;
			51545: outdata = 32'd13991;
			51546: outdata = 32'd13990;
			51547: outdata = 32'd13989;
			51548: outdata = 32'd13988;
			51549: outdata = 32'd13987;
			51550: outdata = 32'd13986;
			51551: outdata = 32'd13985;
			51552: outdata = 32'd13984;
			51553: outdata = 32'd13983;
			51554: outdata = 32'd13982;
			51555: outdata = 32'd13981;
			51556: outdata = 32'd13980;
			51557: outdata = 32'd13979;
			51558: outdata = 32'd13978;
			51559: outdata = 32'd13977;
			51560: outdata = 32'd13976;
			51561: outdata = 32'd13975;
			51562: outdata = 32'd13974;
			51563: outdata = 32'd13973;
			51564: outdata = 32'd13972;
			51565: outdata = 32'd13971;
			51566: outdata = 32'd13970;
			51567: outdata = 32'd13969;
			51568: outdata = 32'd13968;
			51569: outdata = 32'd13967;
			51570: outdata = 32'd13966;
			51571: outdata = 32'd13965;
			51572: outdata = 32'd13964;
			51573: outdata = 32'd13963;
			51574: outdata = 32'd13962;
			51575: outdata = 32'd13961;
			51576: outdata = 32'd13960;
			51577: outdata = 32'd13959;
			51578: outdata = 32'd13958;
			51579: outdata = 32'd13957;
			51580: outdata = 32'd13956;
			51581: outdata = 32'd13955;
			51582: outdata = 32'd13954;
			51583: outdata = 32'd13953;
			51584: outdata = 32'd13952;
			51585: outdata = 32'd13951;
			51586: outdata = 32'd13950;
			51587: outdata = 32'd13949;
			51588: outdata = 32'd13948;
			51589: outdata = 32'd13947;
			51590: outdata = 32'd13946;
			51591: outdata = 32'd13945;
			51592: outdata = 32'd13944;
			51593: outdata = 32'd13943;
			51594: outdata = 32'd13942;
			51595: outdata = 32'd13941;
			51596: outdata = 32'd13940;
			51597: outdata = 32'd13939;
			51598: outdata = 32'd13938;
			51599: outdata = 32'd13937;
			51600: outdata = 32'd13936;
			51601: outdata = 32'd13935;
			51602: outdata = 32'd13934;
			51603: outdata = 32'd13933;
			51604: outdata = 32'd13932;
			51605: outdata = 32'd13931;
			51606: outdata = 32'd13930;
			51607: outdata = 32'd13929;
			51608: outdata = 32'd13928;
			51609: outdata = 32'd13927;
			51610: outdata = 32'd13926;
			51611: outdata = 32'd13925;
			51612: outdata = 32'd13924;
			51613: outdata = 32'd13923;
			51614: outdata = 32'd13922;
			51615: outdata = 32'd13921;
			51616: outdata = 32'd13920;
			51617: outdata = 32'd13919;
			51618: outdata = 32'd13918;
			51619: outdata = 32'd13917;
			51620: outdata = 32'd13916;
			51621: outdata = 32'd13915;
			51622: outdata = 32'd13914;
			51623: outdata = 32'd13913;
			51624: outdata = 32'd13912;
			51625: outdata = 32'd13911;
			51626: outdata = 32'd13910;
			51627: outdata = 32'd13909;
			51628: outdata = 32'd13908;
			51629: outdata = 32'd13907;
			51630: outdata = 32'd13906;
			51631: outdata = 32'd13905;
			51632: outdata = 32'd13904;
			51633: outdata = 32'd13903;
			51634: outdata = 32'd13902;
			51635: outdata = 32'd13901;
			51636: outdata = 32'd13900;
			51637: outdata = 32'd13899;
			51638: outdata = 32'd13898;
			51639: outdata = 32'd13897;
			51640: outdata = 32'd13896;
			51641: outdata = 32'd13895;
			51642: outdata = 32'd13894;
			51643: outdata = 32'd13893;
			51644: outdata = 32'd13892;
			51645: outdata = 32'd13891;
			51646: outdata = 32'd13890;
			51647: outdata = 32'd13889;
			51648: outdata = 32'd13888;
			51649: outdata = 32'd13887;
			51650: outdata = 32'd13886;
			51651: outdata = 32'd13885;
			51652: outdata = 32'd13884;
			51653: outdata = 32'd13883;
			51654: outdata = 32'd13882;
			51655: outdata = 32'd13881;
			51656: outdata = 32'd13880;
			51657: outdata = 32'd13879;
			51658: outdata = 32'd13878;
			51659: outdata = 32'd13877;
			51660: outdata = 32'd13876;
			51661: outdata = 32'd13875;
			51662: outdata = 32'd13874;
			51663: outdata = 32'd13873;
			51664: outdata = 32'd13872;
			51665: outdata = 32'd13871;
			51666: outdata = 32'd13870;
			51667: outdata = 32'd13869;
			51668: outdata = 32'd13868;
			51669: outdata = 32'd13867;
			51670: outdata = 32'd13866;
			51671: outdata = 32'd13865;
			51672: outdata = 32'd13864;
			51673: outdata = 32'd13863;
			51674: outdata = 32'd13862;
			51675: outdata = 32'd13861;
			51676: outdata = 32'd13860;
			51677: outdata = 32'd13859;
			51678: outdata = 32'd13858;
			51679: outdata = 32'd13857;
			51680: outdata = 32'd13856;
			51681: outdata = 32'd13855;
			51682: outdata = 32'd13854;
			51683: outdata = 32'd13853;
			51684: outdata = 32'd13852;
			51685: outdata = 32'd13851;
			51686: outdata = 32'd13850;
			51687: outdata = 32'd13849;
			51688: outdata = 32'd13848;
			51689: outdata = 32'd13847;
			51690: outdata = 32'd13846;
			51691: outdata = 32'd13845;
			51692: outdata = 32'd13844;
			51693: outdata = 32'd13843;
			51694: outdata = 32'd13842;
			51695: outdata = 32'd13841;
			51696: outdata = 32'd13840;
			51697: outdata = 32'd13839;
			51698: outdata = 32'd13838;
			51699: outdata = 32'd13837;
			51700: outdata = 32'd13836;
			51701: outdata = 32'd13835;
			51702: outdata = 32'd13834;
			51703: outdata = 32'd13833;
			51704: outdata = 32'd13832;
			51705: outdata = 32'd13831;
			51706: outdata = 32'd13830;
			51707: outdata = 32'd13829;
			51708: outdata = 32'd13828;
			51709: outdata = 32'd13827;
			51710: outdata = 32'd13826;
			51711: outdata = 32'd13825;
			51712: outdata = 32'd13824;
			51713: outdata = 32'd13823;
			51714: outdata = 32'd13822;
			51715: outdata = 32'd13821;
			51716: outdata = 32'd13820;
			51717: outdata = 32'd13819;
			51718: outdata = 32'd13818;
			51719: outdata = 32'd13817;
			51720: outdata = 32'd13816;
			51721: outdata = 32'd13815;
			51722: outdata = 32'd13814;
			51723: outdata = 32'd13813;
			51724: outdata = 32'd13812;
			51725: outdata = 32'd13811;
			51726: outdata = 32'd13810;
			51727: outdata = 32'd13809;
			51728: outdata = 32'd13808;
			51729: outdata = 32'd13807;
			51730: outdata = 32'd13806;
			51731: outdata = 32'd13805;
			51732: outdata = 32'd13804;
			51733: outdata = 32'd13803;
			51734: outdata = 32'd13802;
			51735: outdata = 32'd13801;
			51736: outdata = 32'd13800;
			51737: outdata = 32'd13799;
			51738: outdata = 32'd13798;
			51739: outdata = 32'd13797;
			51740: outdata = 32'd13796;
			51741: outdata = 32'd13795;
			51742: outdata = 32'd13794;
			51743: outdata = 32'd13793;
			51744: outdata = 32'd13792;
			51745: outdata = 32'd13791;
			51746: outdata = 32'd13790;
			51747: outdata = 32'd13789;
			51748: outdata = 32'd13788;
			51749: outdata = 32'd13787;
			51750: outdata = 32'd13786;
			51751: outdata = 32'd13785;
			51752: outdata = 32'd13784;
			51753: outdata = 32'd13783;
			51754: outdata = 32'd13782;
			51755: outdata = 32'd13781;
			51756: outdata = 32'd13780;
			51757: outdata = 32'd13779;
			51758: outdata = 32'd13778;
			51759: outdata = 32'd13777;
			51760: outdata = 32'd13776;
			51761: outdata = 32'd13775;
			51762: outdata = 32'd13774;
			51763: outdata = 32'd13773;
			51764: outdata = 32'd13772;
			51765: outdata = 32'd13771;
			51766: outdata = 32'd13770;
			51767: outdata = 32'd13769;
			51768: outdata = 32'd13768;
			51769: outdata = 32'd13767;
			51770: outdata = 32'd13766;
			51771: outdata = 32'd13765;
			51772: outdata = 32'd13764;
			51773: outdata = 32'd13763;
			51774: outdata = 32'd13762;
			51775: outdata = 32'd13761;
			51776: outdata = 32'd13760;
			51777: outdata = 32'd13759;
			51778: outdata = 32'd13758;
			51779: outdata = 32'd13757;
			51780: outdata = 32'd13756;
			51781: outdata = 32'd13755;
			51782: outdata = 32'd13754;
			51783: outdata = 32'd13753;
			51784: outdata = 32'd13752;
			51785: outdata = 32'd13751;
			51786: outdata = 32'd13750;
			51787: outdata = 32'd13749;
			51788: outdata = 32'd13748;
			51789: outdata = 32'd13747;
			51790: outdata = 32'd13746;
			51791: outdata = 32'd13745;
			51792: outdata = 32'd13744;
			51793: outdata = 32'd13743;
			51794: outdata = 32'd13742;
			51795: outdata = 32'd13741;
			51796: outdata = 32'd13740;
			51797: outdata = 32'd13739;
			51798: outdata = 32'd13738;
			51799: outdata = 32'd13737;
			51800: outdata = 32'd13736;
			51801: outdata = 32'd13735;
			51802: outdata = 32'd13734;
			51803: outdata = 32'd13733;
			51804: outdata = 32'd13732;
			51805: outdata = 32'd13731;
			51806: outdata = 32'd13730;
			51807: outdata = 32'd13729;
			51808: outdata = 32'd13728;
			51809: outdata = 32'd13727;
			51810: outdata = 32'd13726;
			51811: outdata = 32'd13725;
			51812: outdata = 32'd13724;
			51813: outdata = 32'd13723;
			51814: outdata = 32'd13722;
			51815: outdata = 32'd13721;
			51816: outdata = 32'd13720;
			51817: outdata = 32'd13719;
			51818: outdata = 32'd13718;
			51819: outdata = 32'd13717;
			51820: outdata = 32'd13716;
			51821: outdata = 32'd13715;
			51822: outdata = 32'd13714;
			51823: outdata = 32'd13713;
			51824: outdata = 32'd13712;
			51825: outdata = 32'd13711;
			51826: outdata = 32'd13710;
			51827: outdata = 32'd13709;
			51828: outdata = 32'd13708;
			51829: outdata = 32'd13707;
			51830: outdata = 32'd13706;
			51831: outdata = 32'd13705;
			51832: outdata = 32'd13704;
			51833: outdata = 32'd13703;
			51834: outdata = 32'd13702;
			51835: outdata = 32'd13701;
			51836: outdata = 32'd13700;
			51837: outdata = 32'd13699;
			51838: outdata = 32'd13698;
			51839: outdata = 32'd13697;
			51840: outdata = 32'd13696;
			51841: outdata = 32'd13695;
			51842: outdata = 32'd13694;
			51843: outdata = 32'd13693;
			51844: outdata = 32'd13692;
			51845: outdata = 32'd13691;
			51846: outdata = 32'd13690;
			51847: outdata = 32'd13689;
			51848: outdata = 32'd13688;
			51849: outdata = 32'd13687;
			51850: outdata = 32'd13686;
			51851: outdata = 32'd13685;
			51852: outdata = 32'd13684;
			51853: outdata = 32'd13683;
			51854: outdata = 32'd13682;
			51855: outdata = 32'd13681;
			51856: outdata = 32'd13680;
			51857: outdata = 32'd13679;
			51858: outdata = 32'd13678;
			51859: outdata = 32'd13677;
			51860: outdata = 32'd13676;
			51861: outdata = 32'd13675;
			51862: outdata = 32'd13674;
			51863: outdata = 32'd13673;
			51864: outdata = 32'd13672;
			51865: outdata = 32'd13671;
			51866: outdata = 32'd13670;
			51867: outdata = 32'd13669;
			51868: outdata = 32'd13668;
			51869: outdata = 32'd13667;
			51870: outdata = 32'd13666;
			51871: outdata = 32'd13665;
			51872: outdata = 32'd13664;
			51873: outdata = 32'd13663;
			51874: outdata = 32'd13662;
			51875: outdata = 32'd13661;
			51876: outdata = 32'd13660;
			51877: outdata = 32'd13659;
			51878: outdata = 32'd13658;
			51879: outdata = 32'd13657;
			51880: outdata = 32'd13656;
			51881: outdata = 32'd13655;
			51882: outdata = 32'd13654;
			51883: outdata = 32'd13653;
			51884: outdata = 32'd13652;
			51885: outdata = 32'd13651;
			51886: outdata = 32'd13650;
			51887: outdata = 32'd13649;
			51888: outdata = 32'd13648;
			51889: outdata = 32'd13647;
			51890: outdata = 32'd13646;
			51891: outdata = 32'd13645;
			51892: outdata = 32'd13644;
			51893: outdata = 32'd13643;
			51894: outdata = 32'd13642;
			51895: outdata = 32'd13641;
			51896: outdata = 32'd13640;
			51897: outdata = 32'd13639;
			51898: outdata = 32'd13638;
			51899: outdata = 32'd13637;
			51900: outdata = 32'd13636;
			51901: outdata = 32'd13635;
			51902: outdata = 32'd13634;
			51903: outdata = 32'd13633;
			51904: outdata = 32'd13632;
			51905: outdata = 32'd13631;
			51906: outdata = 32'd13630;
			51907: outdata = 32'd13629;
			51908: outdata = 32'd13628;
			51909: outdata = 32'd13627;
			51910: outdata = 32'd13626;
			51911: outdata = 32'd13625;
			51912: outdata = 32'd13624;
			51913: outdata = 32'd13623;
			51914: outdata = 32'd13622;
			51915: outdata = 32'd13621;
			51916: outdata = 32'd13620;
			51917: outdata = 32'd13619;
			51918: outdata = 32'd13618;
			51919: outdata = 32'd13617;
			51920: outdata = 32'd13616;
			51921: outdata = 32'd13615;
			51922: outdata = 32'd13614;
			51923: outdata = 32'd13613;
			51924: outdata = 32'd13612;
			51925: outdata = 32'd13611;
			51926: outdata = 32'd13610;
			51927: outdata = 32'd13609;
			51928: outdata = 32'd13608;
			51929: outdata = 32'd13607;
			51930: outdata = 32'd13606;
			51931: outdata = 32'd13605;
			51932: outdata = 32'd13604;
			51933: outdata = 32'd13603;
			51934: outdata = 32'd13602;
			51935: outdata = 32'd13601;
			51936: outdata = 32'd13600;
			51937: outdata = 32'd13599;
			51938: outdata = 32'd13598;
			51939: outdata = 32'd13597;
			51940: outdata = 32'd13596;
			51941: outdata = 32'd13595;
			51942: outdata = 32'd13594;
			51943: outdata = 32'd13593;
			51944: outdata = 32'd13592;
			51945: outdata = 32'd13591;
			51946: outdata = 32'd13590;
			51947: outdata = 32'd13589;
			51948: outdata = 32'd13588;
			51949: outdata = 32'd13587;
			51950: outdata = 32'd13586;
			51951: outdata = 32'd13585;
			51952: outdata = 32'd13584;
			51953: outdata = 32'd13583;
			51954: outdata = 32'd13582;
			51955: outdata = 32'd13581;
			51956: outdata = 32'd13580;
			51957: outdata = 32'd13579;
			51958: outdata = 32'd13578;
			51959: outdata = 32'd13577;
			51960: outdata = 32'd13576;
			51961: outdata = 32'd13575;
			51962: outdata = 32'd13574;
			51963: outdata = 32'd13573;
			51964: outdata = 32'd13572;
			51965: outdata = 32'd13571;
			51966: outdata = 32'd13570;
			51967: outdata = 32'd13569;
			51968: outdata = 32'd13568;
			51969: outdata = 32'd13567;
			51970: outdata = 32'd13566;
			51971: outdata = 32'd13565;
			51972: outdata = 32'd13564;
			51973: outdata = 32'd13563;
			51974: outdata = 32'd13562;
			51975: outdata = 32'd13561;
			51976: outdata = 32'd13560;
			51977: outdata = 32'd13559;
			51978: outdata = 32'd13558;
			51979: outdata = 32'd13557;
			51980: outdata = 32'd13556;
			51981: outdata = 32'd13555;
			51982: outdata = 32'd13554;
			51983: outdata = 32'd13553;
			51984: outdata = 32'd13552;
			51985: outdata = 32'd13551;
			51986: outdata = 32'd13550;
			51987: outdata = 32'd13549;
			51988: outdata = 32'd13548;
			51989: outdata = 32'd13547;
			51990: outdata = 32'd13546;
			51991: outdata = 32'd13545;
			51992: outdata = 32'd13544;
			51993: outdata = 32'd13543;
			51994: outdata = 32'd13542;
			51995: outdata = 32'd13541;
			51996: outdata = 32'd13540;
			51997: outdata = 32'd13539;
			51998: outdata = 32'd13538;
			51999: outdata = 32'd13537;
			52000: outdata = 32'd13536;
			52001: outdata = 32'd13535;
			52002: outdata = 32'd13534;
			52003: outdata = 32'd13533;
			52004: outdata = 32'd13532;
			52005: outdata = 32'd13531;
			52006: outdata = 32'd13530;
			52007: outdata = 32'd13529;
			52008: outdata = 32'd13528;
			52009: outdata = 32'd13527;
			52010: outdata = 32'd13526;
			52011: outdata = 32'd13525;
			52012: outdata = 32'd13524;
			52013: outdata = 32'd13523;
			52014: outdata = 32'd13522;
			52015: outdata = 32'd13521;
			52016: outdata = 32'd13520;
			52017: outdata = 32'd13519;
			52018: outdata = 32'd13518;
			52019: outdata = 32'd13517;
			52020: outdata = 32'd13516;
			52021: outdata = 32'd13515;
			52022: outdata = 32'd13514;
			52023: outdata = 32'd13513;
			52024: outdata = 32'd13512;
			52025: outdata = 32'd13511;
			52026: outdata = 32'd13510;
			52027: outdata = 32'd13509;
			52028: outdata = 32'd13508;
			52029: outdata = 32'd13507;
			52030: outdata = 32'd13506;
			52031: outdata = 32'd13505;
			52032: outdata = 32'd13504;
			52033: outdata = 32'd13503;
			52034: outdata = 32'd13502;
			52035: outdata = 32'd13501;
			52036: outdata = 32'd13500;
			52037: outdata = 32'd13499;
			52038: outdata = 32'd13498;
			52039: outdata = 32'd13497;
			52040: outdata = 32'd13496;
			52041: outdata = 32'd13495;
			52042: outdata = 32'd13494;
			52043: outdata = 32'd13493;
			52044: outdata = 32'd13492;
			52045: outdata = 32'd13491;
			52046: outdata = 32'd13490;
			52047: outdata = 32'd13489;
			52048: outdata = 32'd13488;
			52049: outdata = 32'd13487;
			52050: outdata = 32'd13486;
			52051: outdata = 32'd13485;
			52052: outdata = 32'd13484;
			52053: outdata = 32'd13483;
			52054: outdata = 32'd13482;
			52055: outdata = 32'd13481;
			52056: outdata = 32'd13480;
			52057: outdata = 32'd13479;
			52058: outdata = 32'd13478;
			52059: outdata = 32'd13477;
			52060: outdata = 32'd13476;
			52061: outdata = 32'd13475;
			52062: outdata = 32'd13474;
			52063: outdata = 32'd13473;
			52064: outdata = 32'd13472;
			52065: outdata = 32'd13471;
			52066: outdata = 32'd13470;
			52067: outdata = 32'd13469;
			52068: outdata = 32'd13468;
			52069: outdata = 32'd13467;
			52070: outdata = 32'd13466;
			52071: outdata = 32'd13465;
			52072: outdata = 32'd13464;
			52073: outdata = 32'd13463;
			52074: outdata = 32'd13462;
			52075: outdata = 32'd13461;
			52076: outdata = 32'd13460;
			52077: outdata = 32'd13459;
			52078: outdata = 32'd13458;
			52079: outdata = 32'd13457;
			52080: outdata = 32'd13456;
			52081: outdata = 32'd13455;
			52082: outdata = 32'd13454;
			52083: outdata = 32'd13453;
			52084: outdata = 32'd13452;
			52085: outdata = 32'd13451;
			52086: outdata = 32'd13450;
			52087: outdata = 32'd13449;
			52088: outdata = 32'd13448;
			52089: outdata = 32'd13447;
			52090: outdata = 32'd13446;
			52091: outdata = 32'd13445;
			52092: outdata = 32'd13444;
			52093: outdata = 32'd13443;
			52094: outdata = 32'd13442;
			52095: outdata = 32'd13441;
			52096: outdata = 32'd13440;
			52097: outdata = 32'd13439;
			52098: outdata = 32'd13438;
			52099: outdata = 32'd13437;
			52100: outdata = 32'd13436;
			52101: outdata = 32'd13435;
			52102: outdata = 32'd13434;
			52103: outdata = 32'd13433;
			52104: outdata = 32'd13432;
			52105: outdata = 32'd13431;
			52106: outdata = 32'd13430;
			52107: outdata = 32'd13429;
			52108: outdata = 32'd13428;
			52109: outdata = 32'd13427;
			52110: outdata = 32'd13426;
			52111: outdata = 32'd13425;
			52112: outdata = 32'd13424;
			52113: outdata = 32'd13423;
			52114: outdata = 32'd13422;
			52115: outdata = 32'd13421;
			52116: outdata = 32'd13420;
			52117: outdata = 32'd13419;
			52118: outdata = 32'd13418;
			52119: outdata = 32'd13417;
			52120: outdata = 32'd13416;
			52121: outdata = 32'd13415;
			52122: outdata = 32'd13414;
			52123: outdata = 32'd13413;
			52124: outdata = 32'd13412;
			52125: outdata = 32'd13411;
			52126: outdata = 32'd13410;
			52127: outdata = 32'd13409;
			52128: outdata = 32'd13408;
			52129: outdata = 32'd13407;
			52130: outdata = 32'd13406;
			52131: outdata = 32'd13405;
			52132: outdata = 32'd13404;
			52133: outdata = 32'd13403;
			52134: outdata = 32'd13402;
			52135: outdata = 32'd13401;
			52136: outdata = 32'd13400;
			52137: outdata = 32'd13399;
			52138: outdata = 32'd13398;
			52139: outdata = 32'd13397;
			52140: outdata = 32'd13396;
			52141: outdata = 32'd13395;
			52142: outdata = 32'd13394;
			52143: outdata = 32'd13393;
			52144: outdata = 32'd13392;
			52145: outdata = 32'd13391;
			52146: outdata = 32'd13390;
			52147: outdata = 32'd13389;
			52148: outdata = 32'd13388;
			52149: outdata = 32'd13387;
			52150: outdata = 32'd13386;
			52151: outdata = 32'd13385;
			52152: outdata = 32'd13384;
			52153: outdata = 32'd13383;
			52154: outdata = 32'd13382;
			52155: outdata = 32'd13381;
			52156: outdata = 32'd13380;
			52157: outdata = 32'd13379;
			52158: outdata = 32'd13378;
			52159: outdata = 32'd13377;
			52160: outdata = 32'd13376;
			52161: outdata = 32'd13375;
			52162: outdata = 32'd13374;
			52163: outdata = 32'd13373;
			52164: outdata = 32'd13372;
			52165: outdata = 32'd13371;
			52166: outdata = 32'd13370;
			52167: outdata = 32'd13369;
			52168: outdata = 32'd13368;
			52169: outdata = 32'd13367;
			52170: outdata = 32'd13366;
			52171: outdata = 32'd13365;
			52172: outdata = 32'd13364;
			52173: outdata = 32'd13363;
			52174: outdata = 32'd13362;
			52175: outdata = 32'd13361;
			52176: outdata = 32'd13360;
			52177: outdata = 32'd13359;
			52178: outdata = 32'd13358;
			52179: outdata = 32'd13357;
			52180: outdata = 32'd13356;
			52181: outdata = 32'd13355;
			52182: outdata = 32'd13354;
			52183: outdata = 32'd13353;
			52184: outdata = 32'd13352;
			52185: outdata = 32'd13351;
			52186: outdata = 32'd13350;
			52187: outdata = 32'd13349;
			52188: outdata = 32'd13348;
			52189: outdata = 32'd13347;
			52190: outdata = 32'd13346;
			52191: outdata = 32'd13345;
			52192: outdata = 32'd13344;
			52193: outdata = 32'd13343;
			52194: outdata = 32'd13342;
			52195: outdata = 32'd13341;
			52196: outdata = 32'd13340;
			52197: outdata = 32'd13339;
			52198: outdata = 32'd13338;
			52199: outdata = 32'd13337;
			52200: outdata = 32'd13336;
			52201: outdata = 32'd13335;
			52202: outdata = 32'd13334;
			52203: outdata = 32'd13333;
			52204: outdata = 32'd13332;
			52205: outdata = 32'd13331;
			52206: outdata = 32'd13330;
			52207: outdata = 32'd13329;
			52208: outdata = 32'd13328;
			52209: outdata = 32'd13327;
			52210: outdata = 32'd13326;
			52211: outdata = 32'd13325;
			52212: outdata = 32'd13324;
			52213: outdata = 32'd13323;
			52214: outdata = 32'd13322;
			52215: outdata = 32'd13321;
			52216: outdata = 32'd13320;
			52217: outdata = 32'd13319;
			52218: outdata = 32'd13318;
			52219: outdata = 32'd13317;
			52220: outdata = 32'd13316;
			52221: outdata = 32'd13315;
			52222: outdata = 32'd13314;
			52223: outdata = 32'd13313;
			52224: outdata = 32'd13312;
			52225: outdata = 32'd13311;
			52226: outdata = 32'd13310;
			52227: outdata = 32'd13309;
			52228: outdata = 32'd13308;
			52229: outdata = 32'd13307;
			52230: outdata = 32'd13306;
			52231: outdata = 32'd13305;
			52232: outdata = 32'd13304;
			52233: outdata = 32'd13303;
			52234: outdata = 32'd13302;
			52235: outdata = 32'd13301;
			52236: outdata = 32'd13300;
			52237: outdata = 32'd13299;
			52238: outdata = 32'd13298;
			52239: outdata = 32'd13297;
			52240: outdata = 32'd13296;
			52241: outdata = 32'd13295;
			52242: outdata = 32'd13294;
			52243: outdata = 32'd13293;
			52244: outdata = 32'd13292;
			52245: outdata = 32'd13291;
			52246: outdata = 32'd13290;
			52247: outdata = 32'd13289;
			52248: outdata = 32'd13288;
			52249: outdata = 32'd13287;
			52250: outdata = 32'd13286;
			52251: outdata = 32'd13285;
			52252: outdata = 32'd13284;
			52253: outdata = 32'd13283;
			52254: outdata = 32'd13282;
			52255: outdata = 32'd13281;
			52256: outdata = 32'd13280;
			52257: outdata = 32'd13279;
			52258: outdata = 32'd13278;
			52259: outdata = 32'd13277;
			52260: outdata = 32'd13276;
			52261: outdata = 32'd13275;
			52262: outdata = 32'd13274;
			52263: outdata = 32'd13273;
			52264: outdata = 32'd13272;
			52265: outdata = 32'd13271;
			52266: outdata = 32'd13270;
			52267: outdata = 32'd13269;
			52268: outdata = 32'd13268;
			52269: outdata = 32'd13267;
			52270: outdata = 32'd13266;
			52271: outdata = 32'd13265;
			52272: outdata = 32'd13264;
			52273: outdata = 32'd13263;
			52274: outdata = 32'd13262;
			52275: outdata = 32'd13261;
			52276: outdata = 32'd13260;
			52277: outdata = 32'd13259;
			52278: outdata = 32'd13258;
			52279: outdata = 32'd13257;
			52280: outdata = 32'd13256;
			52281: outdata = 32'd13255;
			52282: outdata = 32'd13254;
			52283: outdata = 32'd13253;
			52284: outdata = 32'd13252;
			52285: outdata = 32'd13251;
			52286: outdata = 32'd13250;
			52287: outdata = 32'd13249;
			52288: outdata = 32'd13248;
			52289: outdata = 32'd13247;
			52290: outdata = 32'd13246;
			52291: outdata = 32'd13245;
			52292: outdata = 32'd13244;
			52293: outdata = 32'd13243;
			52294: outdata = 32'd13242;
			52295: outdata = 32'd13241;
			52296: outdata = 32'd13240;
			52297: outdata = 32'd13239;
			52298: outdata = 32'd13238;
			52299: outdata = 32'd13237;
			52300: outdata = 32'd13236;
			52301: outdata = 32'd13235;
			52302: outdata = 32'd13234;
			52303: outdata = 32'd13233;
			52304: outdata = 32'd13232;
			52305: outdata = 32'd13231;
			52306: outdata = 32'd13230;
			52307: outdata = 32'd13229;
			52308: outdata = 32'd13228;
			52309: outdata = 32'd13227;
			52310: outdata = 32'd13226;
			52311: outdata = 32'd13225;
			52312: outdata = 32'd13224;
			52313: outdata = 32'd13223;
			52314: outdata = 32'd13222;
			52315: outdata = 32'd13221;
			52316: outdata = 32'd13220;
			52317: outdata = 32'd13219;
			52318: outdata = 32'd13218;
			52319: outdata = 32'd13217;
			52320: outdata = 32'd13216;
			52321: outdata = 32'd13215;
			52322: outdata = 32'd13214;
			52323: outdata = 32'd13213;
			52324: outdata = 32'd13212;
			52325: outdata = 32'd13211;
			52326: outdata = 32'd13210;
			52327: outdata = 32'd13209;
			52328: outdata = 32'd13208;
			52329: outdata = 32'd13207;
			52330: outdata = 32'd13206;
			52331: outdata = 32'd13205;
			52332: outdata = 32'd13204;
			52333: outdata = 32'd13203;
			52334: outdata = 32'd13202;
			52335: outdata = 32'd13201;
			52336: outdata = 32'd13200;
			52337: outdata = 32'd13199;
			52338: outdata = 32'd13198;
			52339: outdata = 32'd13197;
			52340: outdata = 32'd13196;
			52341: outdata = 32'd13195;
			52342: outdata = 32'd13194;
			52343: outdata = 32'd13193;
			52344: outdata = 32'd13192;
			52345: outdata = 32'd13191;
			52346: outdata = 32'd13190;
			52347: outdata = 32'd13189;
			52348: outdata = 32'd13188;
			52349: outdata = 32'd13187;
			52350: outdata = 32'd13186;
			52351: outdata = 32'd13185;
			52352: outdata = 32'd13184;
			52353: outdata = 32'd13183;
			52354: outdata = 32'd13182;
			52355: outdata = 32'd13181;
			52356: outdata = 32'd13180;
			52357: outdata = 32'd13179;
			52358: outdata = 32'd13178;
			52359: outdata = 32'd13177;
			52360: outdata = 32'd13176;
			52361: outdata = 32'd13175;
			52362: outdata = 32'd13174;
			52363: outdata = 32'd13173;
			52364: outdata = 32'd13172;
			52365: outdata = 32'd13171;
			52366: outdata = 32'd13170;
			52367: outdata = 32'd13169;
			52368: outdata = 32'd13168;
			52369: outdata = 32'd13167;
			52370: outdata = 32'd13166;
			52371: outdata = 32'd13165;
			52372: outdata = 32'd13164;
			52373: outdata = 32'd13163;
			52374: outdata = 32'd13162;
			52375: outdata = 32'd13161;
			52376: outdata = 32'd13160;
			52377: outdata = 32'd13159;
			52378: outdata = 32'd13158;
			52379: outdata = 32'd13157;
			52380: outdata = 32'd13156;
			52381: outdata = 32'd13155;
			52382: outdata = 32'd13154;
			52383: outdata = 32'd13153;
			52384: outdata = 32'd13152;
			52385: outdata = 32'd13151;
			52386: outdata = 32'd13150;
			52387: outdata = 32'd13149;
			52388: outdata = 32'd13148;
			52389: outdata = 32'd13147;
			52390: outdata = 32'd13146;
			52391: outdata = 32'd13145;
			52392: outdata = 32'd13144;
			52393: outdata = 32'd13143;
			52394: outdata = 32'd13142;
			52395: outdata = 32'd13141;
			52396: outdata = 32'd13140;
			52397: outdata = 32'd13139;
			52398: outdata = 32'd13138;
			52399: outdata = 32'd13137;
			52400: outdata = 32'd13136;
			52401: outdata = 32'd13135;
			52402: outdata = 32'd13134;
			52403: outdata = 32'd13133;
			52404: outdata = 32'd13132;
			52405: outdata = 32'd13131;
			52406: outdata = 32'd13130;
			52407: outdata = 32'd13129;
			52408: outdata = 32'd13128;
			52409: outdata = 32'd13127;
			52410: outdata = 32'd13126;
			52411: outdata = 32'd13125;
			52412: outdata = 32'd13124;
			52413: outdata = 32'd13123;
			52414: outdata = 32'd13122;
			52415: outdata = 32'd13121;
			52416: outdata = 32'd13120;
			52417: outdata = 32'd13119;
			52418: outdata = 32'd13118;
			52419: outdata = 32'd13117;
			52420: outdata = 32'd13116;
			52421: outdata = 32'd13115;
			52422: outdata = 32'd13114;
			52423: outdata = 32'd13113;
			52424: outdata = 32'd13112;
			52425: outdata = 32'd13111;
			52426: outdata = 32'd13110;
			52427: outdata = 32'd13109;
			52428: outdata = 32'd13108;
			52429: outdata = 32'd13107;
			52430: outdata = 32'd13106;
			52431: outdata = 32'd13105;
			52432: outdata = 32'd13104;
			52433: outdata = 32'd13103;
			52434: outdata = 32'd13102;
			52435: outdata = 32'd13101;
			52436: outdata = 32'd13100;
			52437: outdata = 32'd13099;
			52438: outdata = 32'd13098;
			52439: outdata = 32'd13097;
			52440: outdata = 32'd13096;
			52441: outdata = 32'd13095;
			52442: outdata = 32'd13094;
			52443: outdata = 32'd13093;
			52444: outdata = 32'd13092;
			52445: outdata = 32'd13091;
			52446: outdata = 32'd13090;
			52447: outdata = 32'd13089;
			52448: outdata = 32'd13088;
			52449: outdata = 32'd13087;
			52450: outdata = 32'd13086;
			52451: outdata = 32'd13085;
			52452: outdata = 32'd13084;
			52453: outdata = 32'd13083;
			52454: outdata = 32'd13082;
			52455: outdata = 32'd13081;
			52456: outdata = 32'd13080;
			52457: outdata = 32'd13079;
			52458: outdata = 32'd13078;
			52459: outdata = 32'd13077;
			52460: outdata = 32'd13076;
			52461: outdata = 32'd13075;
			52462: outdata = 32'd13074;
			52463: outdata = 32'd13073;
			52464: outdata = 32'd13072;
			52465: outdata = 32'd13071;
			52466: outdata = 32'd13070;
			52467: outdata = 32'd13069;
			52468: outdata = 32'd13068;
			52469: outdata = 32'd13067;
			52470: outdata = 32'd13066;
			52471: outdata = 32'd13065;
			52472: outdata = 32'd13064;
			52473: outdata = 32'd13063;
			52474: outdata = 32'd13062;
			52475: outdata = 32'd13061;
			52476: outdata = 32'd13060;
			52477: outdata = 32'd13059;
			52478: outdata = 32'd13058;
			52479: outdata = 32'd13057;
			52480: outdata = 32'd13056;
			52481: outdata = 32'd13055;
			52482: outdata = 32'd13054;
			52483: outdata = 32'd13053;
			52484: outdata = 32'd13052;
			52485: outdata = 32'd13051;
			52486: outdata = 32'd13050;
			52487: outdata = 32'd13049;
			52488: outdata = 32'd13048;
			52489: outdata = 32'd13047;
			52490: outdata = 32'd13046;
			52491: outdata = 32'd13045;
			52492: outdata = 32'd13044;
			52493: outdata = 32'd13043;
			52494: outdata = 32'd13042;
			52495: outdata = 32'd13041;
			52496: outdata = 32'd13040;
			52497: outdata = 32'd13039;
			52498: outdata = 32'd13038;
			52499: outdata = 32'd13037;
			52500: outdata = 32'd13036;
			52501: outdata = 32'd13035;
			52502: outdata = 32'd13034;
			52503: outdata = 32'd13033;
			52504: outdata = 32'd13032;
			52505: outdata = 32'd13031;
			52506: outdata = 32'd13030;
			52507: outdata = 32'd13029;
			52508: outdata = 32'd13028;
			52509: outdata = 32'd13027;
			52510: outdata = 32'd13026;
			52511: outdata = 32'd13025;
			52512: outdata = 32'd13024;
			52513: outdata = 32'd13023;
			52514: outdata = 32'd13022;
			52515: outdata = 32'd13021;
			52516: outdata = 32'd13020;
			52517: outdata = 32'd13019;
			52518: outdata = 32'd13018;
			52519: outdata = 32'd13017;
			52520: outdata = 32'd13016;
			52521: outdata = 32'd13015;
			52522: outdata = 32'd13014;
			52523: outdata = 32'd13013;
			52524: outdata = 32'd13012;
			52525: outdata = 32'd13011;
			52526: outdata = 32'd13010;
			52527: outdata = 32'd13009;
			52528: outdata = 32'd13008;
			52529: outdata = 32'd13007;
			52530: outdata = 32'd13006;
			52531: outdata = 32'd13005;
			52532: outdata = 32'd13004;
			52533: outdata = 32'd13003;
			52534: outdata = 32'd13002;
			52535: outdata = 32'd13001;
			52536: outdata = 32'd13000;
			52537: outdata = 32'd12999;
			52538: outdata = 32'd12998;
			52539: outdata = 32'd12997;
			52540: outdata = 32'd12996;
			52541: outdata = 32'd12995;
			52542: outdata = 32'd12994;
			52543: outdata = 32'd12993;
			52544: outdata = 32'd12992;
			52545: outdata = 32'd12991;
			52546: outdata = 32'd12990;
			52547: outdata = 32'd12989;
			52548: outdata = 32'd12988;
			52549: outdata = 32'd12987;
			52550: outdata = 32'd12986;
			52551: outdata = 32'd12985;
			52552: outdata = 32'd12984;
			52553: outdata = 32'd12983;
			52554: outdata = 32'd12982;
			52555: outdata = 32'd12981;
			52556: outdata = 32'd12980;
			52557: outdata = 32'd12979;
			52558: outdata = 32'd12978;
			52559: outdata = 32'd12977;
			52560: outdata = 32'd12976;
			52561: outdata = 32'd12975;
			52562: outdata = 32'd12974;
			52563: outdata = 32'd12973;
			52564: outdata = 32'd12972;
			52565: outdata = 32'd12971;
			52566: outdata = 32'd12970;
			52567: outdata = 32'd12969;
			52568: outdata = 32'd12968;
			52569: outdata = 32'd12967;
			52570: outdata = 32'd12966;
			52571: outdata = 32'd12965;
			52572: outdata = 32'd12964;
			52573: outdata = 32'd12963;
			52574: outdata = 32'd12962;
			52575: outdata = 32'd12961;
			52576: outdata = 32'd12960;
			52577: outdata = 32'd12959;
			52578: outdata = 32'd12958;
			52579: outdata = 32'd12957;
			52580: outdata = 32'd12956;
			52581: outdata = 32'd12955;
			52582: outdata = 32'd12954;
			52583: outdata = 32'd12953;
			52584: outdata = 32'd12952;
			52585: outdata = 32'd12951;
			52586: outdata = 32'd12950;
			52587: outdata = 32'd12949;
			52588: outdata = 32'd12948;
			52589: outdata = 32'd12947;
			52590: outdata = 32'd12946;
			52591: outdata = 32'd12945;
			52592: outdata = 32'd12944;
			52593: outdata = 32'd12943;
			52594: outdata = 32'd12942;
			52595: outdata = 32'd12941;
			52596: outdata = 32'd12940;
			52597: outdata = 32'd12939;
			52598: outdata = 32'd12938;
			52599: outdata = 32'd12937;
			52600: outdata = 32'd12936;
			52601: outdata = 32'd12935;
			52602: outdata = 32'd12934;
			52603: outdata = 32'd12933;
			52604: outdata = 32'd12932;
			52605: outdata = 32'd12931;
			52606: outdata = 32'd12930;
			52607: outdata = 32'd12929;
			52608: outdata = 32'd12928;
			52609: outdata = 32'd12927;
			52610: outdata = 32'd12926;
			52611: outdata = 32'd12925;
			52612: outdata = 32'd12924;
			52613: outdata = 32'd12923;
			52614: outdata = 32'd12922;
			52615: outdata = 32'd12921;
			52616: outdata = 32'd12920;
			52617: outdata = 32'd12919;
			52618: outdata = 32'd12918;
			52619: outdata = 32'd12917;
			52620: outdata = 32'd12916;
			52621: outdata = 32'd12915;
			52622: outdata = 32'd12914;
			52623: outdata = 32'd12913;
			52624: outdata = 32'd12912;
			52625: outdata = 32'd12911;
			52626: outdata = 32'd12910;
			52627: outdata = 32'd12909;
			52628: outdata = 32'd12908;
			52629: outdata = 32'd12907;
			52630: outdata = 32'd12906;
			52631: outdata = 32'd12905;
			52632: outdata = 32'd12904;
			52633: outdata = 32'd12903;
			52634: outdata = 32'd12902;
			52635: outdata = 32'd12901;
			52636: outdata = 32'd12900;
			52637: outdata = 32'd12899;
			52638: outdata = 32'd12898;
			52639: outdata = 32'd12897;
			52640: outdata = 32'd12896;
			52641: outdata = 32'd12895;
			52642: outdata = 32'd12894;
			52643: outdata = 32'd12893;
			52644: outdata = 32'd12892;
			52645: outdata = 32'd12891;
			52646: outdata = 32'd12890;
			52647: outdata = 32'd12889;
			52648: outdata = 32'd12888;
			52649: outdata = 32'd12887;
			52650: outdata = 32'd12886;
			52651: outdata = 32'd12885;
			52652: outdata = 32'd12884;
			52653: outdata = 32'd12883;
			52654: outdata = 32'd12882;
			52655: outdata = 32'd12881;
			52656: outdata = 32'd12880;
			52657: outdata = 32'd12879;
			52658: outdata = 32'd12878;
			52659: outdata = 32'd12877;
			52660: outdata = 32'd12876;
			52661: outdata = 32'd12875;
			52662: outdata = 32'd12874;
			52663: outdata = 32'd12873;
			52664: outdata = 32'd12872;
			52665: outdata = 32'd12871;
			52666: outdata = 32'd12870;
			52667: outdata = 32'd12869;
			52668: outdata = 32'd12868;
			52669: outdata = 32'd12867;
			52670: outdata = 32'd12866;
			52671: outdata = 32'd12865;
			52672: outdata = 32'd12864;
			52673: outdata = 32'd12863;
			52674: outdata = 32'd12862;
			52675: outdata = 32'd12861;
			52676: outdata = 32'd12860;
			52677: outdata = 32'd12859;
			52678: outdata = 32'd12858;
			52679: outdata = 32'd12857;
			52680: outdata = 32'd12856;
			52681: outdata = 32'd12855;
			52682: outdata = 32'd12854;
			52683: outdata = 32'd12853;
			52684: outdata = 32'd12852;
			52685: outdata = 32'd12851;
			52686: outdata = 32'd12850;
			52687: outdata = 32'd12849;
			52688: outdata = 32'd12848;
			52689: outdata = 32'd12847;
			52690: outdata = 32'd12846;
			52691: outdata = 32'd12845;
			52692: outdata = 32'd12844;
			52693: outdata = 32'd12843;
			52694: outdata = 32'd12842;
			52695: outdata = 32'd12841;
			52696: outdata = 32'd12840;
			52697: outdata = 32'd12839;
			52698: outdata = 32'd12838;
			52699: outdata = 32'd12837;
			52700: outdata = 32'd12836;
			52701: outdata = 32'd12835;
			52702: outdata = 32'd12834;
			52703: outdata = 32'd12833;
			52704: outdata = 32'd12832;
			52705: outdata = 32'd12831;
			52706: outdata = 32'd12830;
			52707: outdata = 32'd12829;
			52708: outdata = 32'd12828;
			52709: outdata = 32'd12827;
			52710: outdata = 32'd12826;
			52711: outdata = 32'd12825;
			52712: outdata = 32'd12824;
			52713: outdata = 32'd12823;
			52714: outdata = 32'd12822;
			52715: outdata = 32'd12821;
			52716: outdata = 32'd12820;
			52717: outdata = 32'd12819;
			52718: outdata = 32'd12818;
			52719: outdata = 32'd12817;
			52720: outdata = 32'd12816;
			52721: outdata = 32'd12815;
			52722: outdata = 32'd12814;
			52723: outdata = 32'd12813;
			52724: outdata = 32'd12812;
			52725: outdata = 32'd12811;
			52726: outdata = 32'd12810;
			52727: outdata = 32'd12809;
			52728: outdata = 32'd12808;
			52729: outdata = 32'd12807;
			52730: outdata = 32'd12806;
			52731: outdata = 32'd12805;
			52732: outdata = 32'd12804;
			52733: outdata = 32'd12803;
			52734: outdata = 32'd12802;
			52735: outdata = 32'd12801;
			52736: outdata = 32'd12800;
			52737: outdata = 32'd12799;
			52738: outdata = 32'd12798;
			52739: outdata = 32'd12797;
			52740: outdata = 32'd12796;
			52741: outdata = 32'd12795;
			52742: outdata = 32'd12794;
			52743: outdata = 32'd12793;
			52744: outdata = 32'd12792;
			52745: outdata = 32'd12791;
			52746: outdata = 32'd12790;
			52747: outdata = 32'd12789;
			52748: outdata = 32'd12788;
			52749: outdata = 32'd12787;
			52750: outdata = 32'd12786;
			52751: outdata = 32'd12785;
			52752: outdata = 32'd12784;
			52753: outdata = 32'd12783;
			52754: outdata = 32'd12782;
			52755: outdata = 32'd12781;
			52756: outdata = 32'd12780;
			52757: outdata = 32'd12779;
			52758: outdata = 32'd12778;
			52759: outdata = 32'd12777;
			52760: outdata = 32'd12776;
			52761: outdata = 32'd12775;
			52762: outdata = 32'd12774;
			52763: outdata = 32'd12773;
			52764: outdata = 32'd12772;
			52765: outdata = 32'd12771;
			52766: outdata = 32'd12770;
			52767: outdata = 32'd12769;
			52768: outdata = 32'd12768;
			52769: outdata = 32'd12767;
			52770: outdata = 32'd12766;
			52771: outdata = 32'd12765;
			52772: outdata = 32'd12764;
			52773: outdata = 32'd12763;
			52774: outdata = 32'd12762;
			52775: outdata = 32'd12761;
			52776: outdata = 32'd12760;
			52777: outdata = 32'd12759;
			52778: outdata = 32'd12758;
			52779: outdata = 32'd12757;
			52780: outdata = 32'd12756;
			52781: outdata = 32'd12755;
			52782: outdata = 32'd12754;
			52783: outdata = 32'd12753;
			52784: outdata = 32'd12752;
			52785: outdata = 32'd12751;
			52786: outdata = 32'd12750;
			52787: outdata = 32'd12749;
			52788: outdata = 32'd12748;
			52789: outdata = 32'd12747;
			52790: outdata = 32'd12746;
			52791: outdata = 32'd12745;
			52792: outdata = 32'd12744;
			52793: outdata = 32'd12743;
			52794: outdata = 32'd12742;
			52795: outdata = 32'd12741;
			52796: outdata = 32'd12740;
			52797: outdata = 32'd12739;
			52798: outdata = 32'd12738;
			52799: outdata = 32'd12737;
			52800: outdata = 32'd12736;
			52801: outdata = 32'd12735;
			52802: outdata = 32'd12734;
			52803: outdata = 32'd12733;
			52804: outdata = 32'd12732;
			52805: outdata = 32'd12731;
			52806: outdata = 32'd12730;
			52807: outdata = 32'd12729;
			52808: outdata = 32'd12728;
			52809: outdata = 32'd12727;
			52810: outdata = 32'd12726;
			52811: outdata = 32'd12725;
			52812: outdata = 32'd12724;
			52813: outdata = 32'd12723;
			52814: outdata = 32'd12722;
			52815: outdata = 32'd12721;
			52816: outdata = 32'd12720;
			52817: outdata = 32'd12719;
			52818: outdata = 32'd12718;
			52819: outdata = 32'd12717;
			52820: outdata = 32'd12716;
			52821: outdata = 32'd12715;
			52822: outdata = 32'd12714;
			52823: outdata = 32'd12713;
			52824: outdata = 32'd12712;
			52825: outdata = 32'd12711;
			52826: outdata = 32'd12710;
			52827: outdata = 32'd12709;
			52828: outdata = 32'd12708;
			52829: outdata = 32'd12707;
			52830: outdata = 32'd12706;
			52831: outdata = 32'd12705;
			52832: outdata = 32'd12704;
			52833: outdata = 32'd12703;
			52834: outdata = 32'd12702;
			52835: outdata = 32'd12701;
			52836: outdata = 32'd12700;
			52837: outdata = 32'd12699;
			52838: outdata = 32'd12698;
			52839: outdata = 32'd12697;
			52840: outdata = 32'd12696;
			52841: outdata = 32'd12695;
			52842: outdata = 32'd12694;
			52843: outdata = 32'd12693;
			52844: outdata = 32'd12692;
			52845: outdata = 32'd12691;
			52846: outdata = 32'd12690;
			52847: outdata = 32'd12689;
			52848: outdata = 32'd12688;
			52849: outdata = 32'd12687;
			52850: outdata = 32'd12686;
			52851: outdata = 32'd12685;
			52852: outdata = 32'd12684;
			52853: outdata = 32'd12683;
			52854: outdata = 32'd12682;
			52855: outdata = 32'd12681;
			52856: outdata = 32'd12680;
			52857: outdata = 32'd12679;
			52858: outdata = 32'd12678;
			52859: outdata = 32'd12677;
			52860: outdata = 32'd12676;
			52861: outdata = 32'd12675;
			52862: outdata = 32'd12674;
			52863: outdata = 32'd12673;
			52864: outdata = 32'd12672;
			52865: outdata = 32'd12671;
			52866: outdata = 32'd12670;
			52867: outdata = 32'd12669;
			52868: outdata = 32'd12668;
			52869: outdata = 32'd12667;
			52870: outdata = 32'd12666;
			52871: outdata = 32'd12665;
			52872: outdata = 32'd12664;
			52873: outdata = 32'd12663;
			52874: outdata = 32'd12662;
			52875: outdata = 32'd12661;
			52876: outdata = 32'd12660;
			52877: outdata = 32'd12659;
			52878: outdata = 32'd12658;
			52879: outdata = 32'd12657;
			52880: outdata = 32'd12656;
			52881: outdata = 32'd12655;
			52882: outdata = 32'd12654;
			52883: outdata = 32'd12653;
			52884: outdata = 32'd12652;
			52885: outdata = 32'd12651;
			52886: outdata = 32'd12650;
			52887: outdata = 32'd12649;
			52888: outdata = 32'd12648;
			52889: outdata = 32'd12647;
			52890: outdata = 32'd12646;
			52891: outdata = 32'd12645;
			52892: outdata = 32'd12644;
			52893: outdata = 32'd12643;
			52894: outdata = 32'd12642;
			52895: outdata = 32'd12641;
			52896: outdata = 32'd12640;
			52897: outdata = 32'd12639;
			52898: outdata = 32'd12638;
			52899: outdata = 32'd12637;
			52900: outdata = 32'd12636;
			52901: outdata = 32'd12635;
			52902: outdata = 32'd12634;
			52903: outdata = 32'd12633;
			52904: outdata = 32'd12632;
			52905: outdata = 32'd12631;
			52906: outdata = 32'd12630;
			52907: outdata = 32'd12629;
			52908: outdata = 32'd12628;
			52909: outdata = 32'd12627;
			52910: outdata = 32'd12626;
			52911: outdata = 32'd12625;
			52912: outdata = 32'd12624;
			52913: outdata = 32'd12623;
			52914: outdata = 32'd12622;
			52915: outdata = 32'd12621;
			52916: outdata = 32'd12620;
			52917: outdata = 32'd12619;
			52918: outdata = 32'd12618;
			52919: outdata = 32'd12617;
			52920: outdata = 32'd12616;
			52921: outdata = 32'd12615;
			52922: outdata = 32'd12614;
			52923: outdata = 32'd12613;
			52924: outdata = 32'd12612;
			52925: outdata = 32'd12611;
			52926: outdata = 32'd12610;
			52927: outdata = 32'd12609;
			52928: outdata = 32'd12608;
			52929: outdata = 32'd12607;
			52930: outdata = 32'd12606;
			52931: outdata = 32'd12605;
			52932: outdata = 32'd12604;
			52933: outdata = 32'd12603;
			52934: outdata = 32'd12602;
			52935: outdata = 32'd12601;
			52936: outdata = 32'd12600;
			52937: outdata = 32'd12599;
			52938: outdata = 32'd12598;
			52939: outdata = 32'd12597;
			52940: outdata = 32'd12596;
			52941: outdata = 32'd12595;
			52942: outdata = 32'd12594;
			52943: outdata = 32'd12593;
			52944: outdata = 32'd12592;
			52945: outdata = 32'd12591;
			52946: outdata = 32'd12590;
			52947: outdata = 32'd12589;
			52948: outdata = 32'd12588;
			52949: outdata = 32'd12587;
			52950: outdata = 32'd12586;
			52951: outdata = 32'd12585;
			52952: outdata = 32'd12584;
			52953: outdata = 32'd12583;
			52954: outdata = 32'd12582;
			52955: outdata = 32'd12581;
			52956: outdata = 32'd12580;
			52957: outdata = 32'd12579;
			52958: outdata = 32'd12578;
			52959: outdata = 32'd12577;
			52960: outdata = 32'd12576;
			52961: outdata = 32'd12575;
			52962: outdata = 32'd12574;
			52963: outdata = 32'd12573;
			52964: outdata = 32'd12572;
			52965: outdata = 32'd12571;
			52966: outdata = 32'd12570;
			52967: outdata = 32'd12569;
			52968: outdata = 32'd12568;
			52969: outdata = 32'd12567;
			52970: outdata = 32'd12566;
			52971: outdata = 32'd12565;
			52972: outdata = 32'd12564;
			52973: outdata = 32'd12563;
			52974: outdata = 32'd12562;
			52975: outdata = 32'd12561;
			52976: outdata = 32'd12560;
			52977: outdata = 32'd12559;
			52978: outdata = 32'd12558;
			52979: outdata = 32'd12557;
			52980: outdata = 32'd12556;
			52981: outdata = 32'd12555;
			52982: outdata = 32'd12554;
			52983: outdata = 32'd12553;
			52984: outdata = 32'd12552;
			52985: outdata = 32'd12551;
			52986: outdata = 32'd12550;
			52987: outdata = 32'd12549;
			52988: outdata = 32'd12548;
			52989: outdata = 32'd12547;
			52990: outdata = 32'd12546;
			52991: outdata = 32'd12545;
			52992: outdata = 32'd12544;
			52993: outdata = 32'd12543;
			52994: outdata = 32'd12542;
			52995: outdata = 32'd12541;
			52996: outdata = 32'd12540;
			52997: outdata = 32'd12539;
			52998: outdata = 32'd12538;
			52999: outdata = 32'd12537;
			53000: outdata = 32'd12536;
			53001: outdata = 32'd12535;
			53002: outdata = 32'd12534;
			53003: outdata = 32'd12533;
			53004: outdata = 32'd12532;
			53005: outdata = 32'd12531;
			53006: outdata = 32'd12530;
			53007: outdata = 32'd12529;
			53008: outdata = 32'd12528;
			53009: outdata = 32'd12527;
			53010: outdata = 32'd12526;
			53011: outdata = 32'd12525;
			53012: outdata = 32'd12524;
			53013: outdata = 32'd12523;
			53014: outdata = 32'd12522;
			53015: outdata = 32'd12521;
			53016: outdata = 32'd12520;
			53017: outdata = 32'd12519;
			53018: outdata = 32'd12518;
			53019: outdata = 32'd12517;
			53020: outdata = 32'd12516;
			53021: outdata = 32'd12515;
			53022: outdata = 32'd12514;
			53023: outdata = 32'd12513;
			53024: outdata = 32'd12512;
			53025: outdata = 32'd12511;
			53026: outdata = 32'd12510;
			53027: outdata = 32'd12509;
			53028: outdata = 32'd12508;
			53029: outdata = 32'd12507;
			53030: outdata = 32'd12506;
			53031: outdata = 32'd12505;
			53032: outdata = 32'd12504;
			53033: outdata = 32'd12503;
			53034: outdata = 32'd12502;
			53035: outdata = 32'd12501;
			53036: outdata = 32'd12500;
			53037: outdata = 32'd12499;
			53038: outdata = 32'd12498;
			53039: outdata = 32'd12497;
			53040: outdata = 32'd12496;
			53041: outdata = 32'd12495;
			53042: outdata = 32'd12494;
			53043: outdata = 32'd12493;
			53044: outdata = 32'd12492;
			53045: outdata = 32'd12491;
			53046: outdata = 32'd12490;
			53047: outdata = 32'd12489;
			53048: outdata = 32'd12488;
			53049: outdata = 32'd12487;
			53050: outdata = 32'd12486;
			53051: outdata = 32'd12485;
			53052: outdata = 32'd12484;
			53053: outdata = 32'd12483;
			53054: outdata = 32'd12482;
			53055: outdata = 32'd12481;
			53056: outdata = 32'd12480;
			53057: outdata = 32'd12479;
			53058: outdata = 32'd12478;
			53059: outdata = 32'd12477;
			53060: outdata = 32'd12476;
			53061: outdata = 32'd12475;
			53062: outdata = 32'd12474;
			53063: outdata = 32'd12473;
			53064: outdata = 32'd12472;
			53065: outdata = 32'd12471;
			53066: outdata = 32'd12470;
			53067: outdata = 32'd12469;
			53068: outdata = 32'd12468;
			53069: outdata = 32'd12467;
			53070: outdata = 32'd12466;
			53071: outdata = 32'd12465;
			53072: outdata = 32'd12464;
			53073: outdata = 32'd12463;
			53074: outdata = 32'd12462;
			53075: outdata = 32'd12461;
			53076: outdata = 32'd12460;
			53077: outdata = 32'd12459;
			53078: outdata = 32'd12458;
			53079: outdata = 32'd12457;
			53080: outdata = 32'd12456;
			53081: outdata = 32'd12455;
			53082: outdata = 32'd12454;
			53083: outdata = 32'd12453;
			53084: outdata = 32'd12452;
			53085: outdata = 32'd12451;
			53086: outdata = 32'd12450;
			53087: outdata = 32'd12449;
			53088: outdata = 32'd12448;
			53089: outdata = 32'd12447;
			53090: outdata = 32'd12446;
			53091: outdata = 32'd12445;
			53092: outdata = 32'd12444;
			53093: outdata = 32'd12443;
			53094: outdata = 32'd12442;
			53095: outdata = 32'd12441;
			53096: outdata = 32'd12440;
			53097: outdata = 32'd12439;
			53098: outdata = 32'd12438;
			53099: outdata = 32'd12437;
			53100: outdata = 32'd12436;
			53101: outdata = 32'd12435;
			53102: outdata = 32'd12434;
			53103: outdata = 32'd12433;
			53104: outdata = 32'd12432;
			53105: outdata = 32'd12431;
			53106: outdata = 32'd12430;
			53107: outdata = 32'd12429;
			53108: outdata = 32'd12428;
			53109: outdata = 32'd12427;
			53110: outdata = 32'd12426;
			53111: outdata = 32'd12425;
			53112: outdata = 32'd12424;
			53113: outdata = 32'd12423;
			53114: outdata = 32'd12422;
			53115: outdata = 32'd12421;
			53116: outdata = 32'd12420;
			53117: outdata = 32'd12419;
			53118: outdata = 32'd12418;
			53119: outdata = 32'd12417;
			53120: outdata = 32'd12416;
			53121: outdata = 32'd12415;
			53122: outdata = 32'd12414;
			53123: outdata = 32'd12413;
			53124: outdata = 32'd12412;
			53125: outdata = 32'd12411;
			53126: outdata = 32'd12410;
			53127: outdata = 32'd12409;
			53128: outdata = 32'd12408;
			53129: outdata = 32'd12407;
			53130: outdata = 32'd12406;
			53131: outdata = 32'd12405;
			53132: outdata = 32'd12404;
			53133: outdata = 32'd12403;
			53134: outdata = 32'd12402;
			53135: outdata = 32'd12401;
			53136: outdata = 32'd12400;
			53137: outdata = 32'd12399;
			53138: outdata = 32'd12398;
			53139: outdata = 32'd12397;
			53140: outdata = 32'd12396;
			53141: outdata = 32'd12395;
			53142: outdata = 32'd12394;
			53143: outdata = 32'd12393;
			53144: outdata = 32'd12392;
			53145: outdata = 32'd12391;
			53146: outdata = 32'd12390;
			53147: outdata = 32'd12389;
			53148: outdata = 32'd12388;
			53149: outdata = 32'd12387;
			53150: outdata = 32'd12386;
			53151: outdata = 32'd12385;
			53152: outdata = 32'd12384;
			53153: outdata = 32'd12383;
			53154: outdata = 32'd12382;
			53155: outdata = 32'd12381;
			53156: outdata = 32'd12380;
			53157: outdata = 32'd12379;
			53158: outdata = 32'd12378;
			53159: outdata = 32'd12377;
			53160: outdata = 32'd12376;
			53161: outdata = 32'd12375;
			53162: outdata = 32'd12374;
			53163: outdata = 32'd12373;
			53164: outdata = 32'd12372;
			53165: outdata = 32'd12371;
			53166: outdata = 32'd12370;
			53167: outdata = 32'd12369;
			53168: outdata = 32'd12368;
			53169: outdata = 32'd12367;
			53170: outdata = 32'd12366;
			53171: outdata = 32'd12365;
			53172: outdata = 32'd12364;
			53173: outdata = 32'd12363;
			53174: outdata = 32'd12362;
			53175: outdata = 32'd12361;
			53176: outdata = 32'd12360;
			53177: outdata = 32'd12359;
			53178: outdata = 32'd12358;
			53179: outdata = 32'd12357;
			53180: outdata = 32'd12356;
			53181: outdata = 32'd12355;
			53182: outdata = 32'd12354;
			53183: outdata = 32'd12353;
			53184: outdata = 32'd12352;
			53185: outdata = 32'd12351;
			53186: outdata = 32'd12350;
			53187: outdata = 32'd12349;
			53188: outdata = 32'd12348;
			53189: outdata = 32'd12347;
			53190: outdata = 32'd12346;
			53191: outdata = 32'd12345;
			53192: outdata = 32'd12344;
			53193: outdata = 32'd12343;
			53194: outdata = 32'd12342;
			53195: outdata = 32'd12341;
			53196: outdata = 32'd12340;
			53197: outdata = 32'd12339;
			53198: outdata = 32'd12338;
			53199: outdata = 32'd12337;
			53200: outdata = 32'd12336;
			53201: outdata = 32'd12335;
			53202: outdata = 32'd12334;
			53203: outdata = 32'd12333;
			53204: outdata = 32'd12332;
			53205: outdata = 32'd12331;
			53206: outdata = 32'd12330;
			53207: outdata = 32'd12329;
			53208: outdata = 32'd12328;
			53209: outdata = 32'd12327;
			53210: outdata = 32'd12326;
			53211: outdata = 32'd12325;
			53212: outdata = 32'd12324;
			53213: outdata = 32'd12323;
			53214: outdata = 32'd12322;
			53215: outdata = 32'd12321;
			53216: outdata = 32'd12320;
			53217: outdata = 32'd12319;
			53218: outdata = 32'd12318;
			53219: outdata = 32'd12317;
			53220: outdata = 32'd12316;
			53221: outdata = 32'd12315;
			53222: outdata = 32'd12314;
			53223: outdata = 32'd12313;
			53224: outdata = 32'd12312;
			53225: outdata = 32'd12311;
			53226: outdata = 32'd12310;
			53227: outdata = 32'd12309;
			53228: outdata = 32'd12308;
			53229: outdata = 32'd12307;
			53230: outdata = 32'd12306;
			53231: outdata = 32'd12305;
			53232: outdata = 32'd12304;
			53233: outdata = 32'd12303;
			53234: outdata = 32'd12302;
			53235: outdata = 32'd12301;
			53236: outdata = 32'd12300;
			53237: outdata = 32'd12299;
			53238: outdata = 32'd12298;
			53239: outdata = 32'd12297;
			53240: outdata = 32'd12296;
			53241: outdata = 32'd12295;
			53242: outdata = 32'd12294;
			53243: outdata = 32'd12293;
			53244: outdata = 32'd12292;
			53245: outdata = 32'd12291;
			53246: outdata = 32'd12290;
			53247: outdata = 32'd12289;
			53248: outdata = 32'd12288;
			53249: outdata = 32'd12287;
			53250: outdata = 32'd12286;
			53251: outdata = 32'd12285;
			53252: outdata = 32'd12284;
			53253: outdata = 32'd12283;
			53254: outdata = 32'd12282;
			53255: outdata = 32'd12281;
			53256: outdata = 32'd12280;
			53257: outdata = 32'd12279;
			53258: outdata = 32'd12278;
			53259: outdata = 32'd12277;
			53260: outdata = 32'd12276;
			53261: outdata = 32'd12275;
			53262: outdata = 32'd12274;
			53263: outdata = 32'd12273;
			53264: outdata = 32'd12272;
			53265: outdata = 32'd12271;
			53266: outdata = 32'd12270;
			53267: outdata = 32'd12269;
			53268: outdata = 32'd12268;
			53269: outdata = 32'd12267;
			53270: outdata = 32'd12266;
			53271: outdata = 32'd12265;
			53272: outdata = 32'd12264;
			53273: outdata = 32'd12263;
			53274: outdata = 32'd12262;
			53275: outdata = 32'd12261;
			53276: outdata = 32'd12260;
			53277: outdata = 32'd12259;
			53278: outdata = 32'd12258;
			53279: outdata = 32'd12257;
			53280: outdata = 32'd12256;
			53281: outdata = 32'd12255;
			53282: outdata = 32'd12254;
			53283: outdata = 32'd12253;
			53284: outdata = 32'd12252;
			53285: outdata = 32'd12251;
			53286: outdata = 32'd12250;
			53287: outdata = 32'd12249;
			53288: outdata = 32'd12248;
			53289: outdata = 32'd12247;
			53290: outdata = 32'd12246;
			53291: outdata = 32'd12245;
			53292: outdata = 32'd12244;
			53293: outdata = 32'd12243;
			53294: outdata = 32'd12242;
			53295: outdata = 32'd12241;
			53296: outdata = 32'd12240;
			53297: outdata = 32'd12239;
			53298: outdata = 32'd12238;
			53299: outdata = 32'd12237;
			53300: outdata = 32'd12236;
			53301: outdata = 32'd12235;
			53302: outdata = 32'd12234;
			53303: outdata = 32'd12233;
			53304: outdata = 32'd12232;
			53305: outdata = 32'd12231;
			53306: outdata = 32'd12230;
			53307: outdata = 32'd12229;
			53308: outdata = 32'd12228;
			53309: outdata = 32'd12227;
			53310: outdata = 32'd12226;
			53311: outdata = 32'd12225;
			53312: outdata = 32'd12224;
			53313: outdata = 32'd12223;
			53314: outdata = 32'd12222;
			53315: outdata = 32'd12221;
			53316: outdata = 32'd12220;
			53317: outdata = 32'd12219;
			53318: outdata = 32'd12218;
			53319: outdata = 32'd12217;
			53320: outdata = 32'd12216;
			53321: outdata = 32'd12215;
			53322: outdata = 32'd12214;
			53323: outdata = 32'd12213;
			53324: outdata = 32'd12212;
			53325: outdata = 32'd12211;
			53326: outdata = 32'd12210;
			53327: outdata = 32'd12209;
			53328: outdata = 32'd12208;
			53329: outdata = 32'd12207;
			53330: outdata = 32'd12206;
			53331: outdata = 32'd12205;
			53332: outdata = 32'd12204;
			53333: outdata = 32'd12203;
			53334: outdata = 32'd12202;
			53335: outdata = 32'd12201;
			53336: outdata = 32'd12200;
			53337: outdata = 32'd12199;
			53338: outdata = 32'd12198;
			53339: outdata = 32'd12197;
			53340: outdata = 32'd12196;
			53341: outdata = 32'd12195;
			53342: outdata = 32'd12194;
			53343: outdata = 32'd12193;
			53344: outdata = 32'd12192;
			53345: outdata = 32'd12191;
			53346: outdata = 32'd12190;
			53347: outdata = 32'd12189;
			53348: outdata = 32'd12188;
			53349: outdata = 32'd12187;
			53350: outdata = 32'd12186;
			53351: outdata = 32'd12185;
			53352: outdata = 32'd12184;
			53353: outdata = 32'd12183;
			53354: outdata = 32'd12182;
			53355: outdata = 32'd12181;
			53356: outdata = 32'd12180;
			53357: outdata = 32'd12179;
			53358: outdata = 32'd12178;
			53359: outdata = 32'd12177;
			53360: outdata = 32'd12176;
			53361: outdata = 32'd12175;
			53362: outdata = 32'd12174;
			53363: outdata = 32'd12173;
			53364: outdata = 32'd12172;
			53365: outdata = 32'd12171;
			53366: outdata = 32'd12170;
			53367: outdata = 32'd12169;
			53368: outdata = 32'd12168;
			53369: outdata = 32'd12167;
			53370: outdata = 32'd12166;
			53371: outdata = 32'd12165;
			53372: outdata = 32'd12164;
			53373: outdata = 32'd12163;
			53374: outdata = 32'd12162;
			53375: outdata = 32'd12161;
			53376: outdata = 32'd12160;
			53377: outdata = 32'd12159;
			53378: outdata = 32'd12158;
			53379: outdata = 32'd12157;
			53380: outdata = 32'd12156;
			53381: outdata = 32'd12155;
			53382: outdata = 32'd12154;
			53383: outdata = 32'd12153;
			53384: outdata = 32'd12152;
			53385: outdata = 32'd12151;
			53386: outdata = 32'd12150;
			53387: outdata = 32'd12149;
			53388: outdata = 32'd12148;
			53389: outdata = 32'd12147;
			53390: outdata = 32'd12146;
			53391: outdata = 32'd12145;
			53392: outdata = 32'd12144;
			53393: outdata = 32'd12143;
			53394: outdata = 32'd12142;
			53395: outdata = 32'd12141;
			53396: outdata = 32'd12140;
			53397: outdata = 32'd12139;
			53398: outdata = 32'd12138;
			53399: outdata = 32'd12137;
			53400: outdata = 32'd12136;
			53401: outdata = 32'd12135;
			53402: outdata = 32'd12134;
			53403: outdata = 32'd12133;
			53404: outdata = 32'd12132;
			53405: outdata = 32'd12131;
			53406: outdata = 32'd12130;
			53407: outdata = 32'd12129;
			53408: outdata = 32'd12128;
			53409: outdata = 32'd12127;
			53410: outdata = 32'd12126;
			53411: outdata = 32'd12125;
			53412: outdata = 32'd12124;
			53413: outdata = 32'd12123;
			53414: outdata = 32'd12122;
			53415: outdata = 32'd12121;
			53416: outdata = 32'd12120;
			53417: outdata = 32'd12119;
			53418: outdata = 32'd12118;
			53419: outdata = 32'd12117;
			53420: outdata = 32'd12116;
			53421: outdata = 32'd12115;
			53422: outdata = 32'd12114;
			53423: outdata = 32'd12113;
			53424: outdata = 32'd12112;
			53425: outdata = 32'd12111;
			53426: outdata = 32'd12110;
			53427: outdata = 32'd12109;
			53428: outdata = 32'd12108;
			53429: outdata = 32'd12107;
			53430: outdata = 32'd12106;
			53431: outdata = 32'd12105;
			53432: outdata = 32'd12104;
			53433: outdata = 32'd12103;
			53434: outdata = 32'd12102;
			53435: outdata = 32'd12101;
			53436: outdata = 32'd12100;
			53437: outdata = 32'd12099;
			53438: outdata = 32'd12098;
			53439: outdata = 32'd12097;
			53440: outdata = 32'd12096;
			53441: outdata = 32'd12095;
			53442: outdata = 32'd12094;
			53443: outdata = 32'd12093;
			53444: outdata = 32'd12092;
			53445: outdata = 32'd12091;
			53446: outdata = 32'd12090;
			53447: outdata = 32'd12089;
			53448: outdata = 32'd12088;
			53449: outdata = 32'd12087;
			53450: outdata = 32'd12086;
			53451: outdata = 32'd12085;
			53452: outdata = 32'd12084;
			53453: outdata = 32'd12083;
			53454: outdata = 32'd12082;
			53455: outdata = 32'd12081;
			53456: outdata = 32'd12080;
			53457: outdata = 32'd12079;
			53458: outdata = 32'd12078;
			53459: outdata = 32'd12077;
			53460: outdata = 32'd12076;
			53461: outdata = 32'd12075;
			53462: outdata = 32'd12074;
			53463: outdata = 32'd12073;
			53464: outdata = 32'd12072;
			53465: outdata = 32'd12071;
			53466: outdata = 32'd12070;
			53467: outdata = 32'd12069;
			53468: outdata = 32'd12068;
			53469: outdata = 32'd12067;
			53470: outdata = 32'd12066;
			53471: outdata = 32'd12065;
			53472: outdata = 32'd12064;
			53473: outdata = 32'd12063;
			53474: outdata = 32'd12062;
			53475: outdata = 32'd12061;
			53476: outdata = 32'd12060;
			53477: outdata = 32'd12059;
			53478: outdata = 32'd12058;
			53479: outdata = 32'd12057;
			53480: outdata = 32'd12056;
			53481: outdata = 32'd12055;
			53482: outdata = 32'd12054;
			53483: outdata = 32'd12053;
			53484: outdata = 32'd12052;
			53485: outdata = 32'd12051;
			53486: outdata = 32'd12050;
			53487: outdata = 32'd12049;
			53488: outdata = 32'd12048;
			53489: outdata = 32'd12047;
			53490: outdata = 32'd12046;
			53491: outdata = 32'd12045;
			53492: outdata = 32'd12044;
			53493: outdata = 32'd12043;
			53494: outdata = 32'd12042;
			53495: outdata = 32'd12041;
			53496: outdata = 32'd12040;
			53497: outdata = 32'd12039;
			53498: outdata = 32'd12038;
			53499: outdata = 32'd12037;
			53500: outdata = 32'd12036;
			53501: outdata = 32'd12035;
			53502: outdata = 32'd12034;
			53503: outdata = 32'd12033;
			53504: outdata = 32'd12032;
			53505: outdata = 32'd12031;
			53506: outdata = 32'd12030;
			53507: outdata = 32'd12029;
			53508: outdata = 32'd12028;
			53509: outdata = 32'd12027;
			53510: outdata = 32'd12026;
			53511: outdata = 32'd12025;
			53512: outdata = 32'd12024;
			53513: outdata = 32'd12023;
			53514: outdata = 32'd12022;
			53515: outdata = 32'd12021;
			53516: outdata = 32'd12020;
			53517: outdata = 32'd12019;
			53518: outdata = 32'd12018;
			53519: outdata = 32'd12017;
			53520: outdata = 32'd12016;
			53521: outdata = 32'd12015;
			53522: outdata = 32'd12014;
			53523: outdata = 32'd12013;
			53524: outdata = 32'd12012;
			53525: outdata = 32'd12011;
			53526: outdata = 32'd12010;
			53527: outdata = 32'd12009;
			53528: outdata = 32'd12008;
			53529: outdata = 32'd12007;
			53530: outdata = 32'd12006;
			53531: outdata = 32'd12005;
			53532: outdata = 32'd12004;
			53533: outdata = 32'd12003;
			53534: outdata = 32'd12002;
			53535: outdata = 32'd12001;
			53536: outdata = 32'd12000;
			53537: outdata = 32'd11999;
			53538: outdata = 32'd11998;
			53539: outdata = 32'd11997;
			53540: outdata = 32'd11996;
			53541: outdata = 32'd11995;
			53542: outdata = 32'd11994;
			53543: outdata = 32'd11993;
			53544: outdata = 32'd11992;
			53545: outdata = 32'd11991;
			53546: outdata = 32'd11990;
			53547: outdata = 32'd11989;
			53548: outdata = 32'd11988;
			53549: outdata = 32'd11987;
			53550: outdata = 32'd11986;
			53551: outdata = 32'd11985;
			53552: outdata = 32'd11984;
			53553: outdata = 32'd11983;
			53554: outdata = 32'd11982;
			53555: outdata = 32'd11981;
			53556: outdata = 32'd11980;
			53557: outdata = 32'd11979;
			53558: outdata = 32'd11978;
			53559: outdata = 32'd11977;
			53560: outdata = 32'd11976;
			53561: outdata = 32'd11975;
			53562: outdata = 32'd11974;
			53563: outdata = 32'd11973;
			53564: outdata = 32'd11972;
			53565: outdata = 32'd11971;
			53566: outdata = 32'd11970;
			53567: outdata = 32'd11969;
			53568: outdata = 32'd11968;
			53569: outdata = 32'd11967;
			53570: outdata = 32'd11966;
			53571: outdata = 32'd11965;
			53572: outdata = 32'd11964;
			53573: outdata = 32'd11963;
			53574: outdata = 32'd11962;
			53575: outdata = 32'd11961;
			53576: outdata = 32'd11960;
			53577: outdata = 32'd11959;
			53578: outdata = 32'd11958;
			53579: outdata = 32'd11957;
			53580: outdata = 32'd11956;
			53581: outdata = 32'd11955;
			53582: outdata = 32'd11954;
			53583: outdata = 32'd11953;
			53584: outdata = 32'd11952;
			53585: outdata = 32'd11951;
			53586: outdata = 32'd11950;
			53587: outdata = 32'd11949;
			53588: outdata = 32'd11948;
			53589: outdata = 32'd11947;
			53590: outdata = 32'd11946;
			53591: outdata = 32'd11945;
			53592: outdata = 32'd11944;
			53593: outdata = 32'd11943;
			53594: outdata = 32'd11942;
			53595: outdata = 32'd11941;
			53596: outdata = 32'd11940;
			53597: outdata = 32'd11939;
			53598: outdata = 32'd11938;
			53599: outdata = 32'd11937;
			53600: outdata = 32'd11936;
			53601: outdata = 32'd11935;
			53602: outdata = 32'd11934;
			53603: outdata = 32'd11933;
			53604: outdata = 32'd11932;
			53605: outdata = 32'd11931;
			53606: outdata = 32'd11930;
			53607: outdata = 32'd11929;
			53608: outdata = 32'd11928;
			53609: outdata = 32'd11927;
			53610: outdata = 32'd11926;
			53611: outdata = 32'd11925;
			53612: outdata = 32'd11924;
			53613: outdata = 32'd11923;
			53614: outdata = 32'd11922;
			53615: outdata = 32'd11921;
			53616: outdata = 32'd11920;
			53617: outdata = 32'd11919;
			53618: outdata = 32'd11918;
			53619: outdata = 32'd11917;
			53620: outdata = 32'd11916;
			53621: outdata = 32'd11915;
			53622: outdata = 32'd11914;
			53623: outdata = 32'd11913;
			53624: outdata = 32'd11912;
			53625: outdata = 32'd11911;
			53626: outdata = 32'd11910;
			53627: outdata = 32'd11909;
			53628: outdata = 32'd11908;
			53629: outdata = 32'd11907;
			53630: outdata = 32'd11906;
			53631: outdata = 32'd11905;
			53632: outdata = 32'd11904;
			53633: outdata = 32'd11903;
			53634: outdata = 32'd11902;
			53635: outdata = 32'd11901;
			53636: outdata = 32'd11900;
			53637: outdata = 32'd11899;
			53638: outdata = 32'd11898;
			53639: outdata = 32'd11897;
			53640: outdata = 32'd11896;
			53641: outdata = 32'd11895;
			53642: outdata = 32'd11894;
			53643: outdata = 32'd11893;
			53644: outdata = 32'd11892;
			53645: outdata = 32'd11891;
			53646: outdata = 32'd11890;
			53647: outdata = 32'd11889;
			53648: outdata = 32'd11888;
			53649: outdata = 32'd11887;
			53650: outdata = 32'd11886;
			53651: outdata = 32'd11885;
			53652: outdata = 32'd11884;
			53653: outdata = 32'd11883;
			53654: outdata = 32'd11882;
			53655: outdata = 32'd11881;
			53656: outdata = 32'd11880;
			53657: outdata = 32'd11879;
			53658: outdata = 32'd11878;
			53659: outdata = 32'd11877;
			53660: outdata = 32'd11876;
			53661: outdata = 32'd11875;
			53662: outdata = 32'd11874;
			53663: outdata = 32'd11873;
			53664: outdata = 32'd11872;
			53665: outdata = 32'd11871;
			53666: outdata = 32'd11870;
			53667: outdata = 32'd11869;
			53668: outdata = 32'd11868;
			53669: outdata = 32'd11867;
			53670: outdata = 32'd11866;
			53671: outdata = 32'd11865;
			53672: outdata = 32'd11864;
			53673: outdata = 32'd11863;
			53674: outdata = 32'd11862;
			53675: outdata = 32'd11861;
			53676: outdata = 32'd11860;
			53677: outdata = 32'd11859;
			53678: outdata = 32'd11858;
			53679: outdata = 32'd11857;
			53680: outdata = 32'd11856;
			53681: outdata = 32'd11855;
			53682: outdata = 32'd11854;
			53683: outdata = 32'd11853;
			53684: outdata = 32'd11852;
			53685: outdata = 32'd11851;
			53686: outdata = 32'd11850;
			53687: outdata = 32'd11849;
			53688: outdata = 32'd11848;
			53689: outdata = 32'd11847;
			53690: outdata = 32'd11846;
			53691: outdata = 32'd11845;
			53692: outdata = 32'd11844;
			53693: outdata = 32'd11843;
			53694: outdata = 32'd11842;
			53695: outdata = 32'd11841;
			53696: outdata = 32'd11840;
			53697: outdata = 32'd11839;
			53698: outdata = 32'd11838;
			53699: outdata = 32'd11837;
			53700: outdata = 32'd11836;
			53701: outdata = 32'd11835;
			53702: outdata = 32'd11834;
			53703: outdata = 32'd11833;
			53704: outdata = 32'd11832;
			53705: outdata = 32'd11831;
			53706: outdata = 32'd11830;
			53707: outdata = 32'd11829;
			53708: outdata = 32'd11828;
			53709: outdata = 32'd11827;
			53710: outdata = 32'd11826;
			53711: outdata = 32'd11825;
			53712: outdata = 32'd11824;
			53713: outdata = 32'd11823;
			53714: outdata = 32'd11822;
			53715: outdata = 32'd11821;
			53716: outdata = 32'd11820;
			53717: outdata = 32'd11819;
			53718: outdata = 32'd11818;
			53719: outdata = 32'd11817;
			53720: outdata = 32'd11816;
			53721: outdata = 32'd11815;
			53722: outdata = 32'd11814;
			53723: outdata = 32'd11813;
			53724: outdata = 32'd11812;
			53725: outdata = 32'd11811;
			53726: outdata = 32'd11810;
			53727: outdata = 32'd11809;
			53728: outdata = 32'd11808;
			53729: outdata = 32'd11807;
			53730: outdata = 32'd11806;
			53731: outdata = 32'd11805;
			53732: outdata = 32'd11804;
			53733: outdata = 32'd11803;
			53734: outdata = 32'd11802;
			53735: outdata = 32'd11801;
			53736: outdata = 32'd11800;
			53737: outdata = 32'd11799;
			53738: outdata = 32'd11798;
			53739: outdata = 32'd11797;
			53740: outdata = 32'd11796;
			53741: outdata = 32'd11795;
			53742: outdata = 32'd11794;
			53743: outdata = 32'd11793;
			53744: outdata = 32'd11792;
			53745: outdata = 32'd11791;
			53746: outdata = 32'd11790;
			53747: outdata = 32'd11789;
			53748: outdata = 32'd11788;
			53749: outdata = 32'd11787;
			53750: outdata = 32'd11786;
			53751: outdata = 32'd11785;
			53752: outdata = 32'd11784;
			53753: outdata = 32'd11783;
			53754: outdata = 32'd11782;
			53755: outdata = 32'd11781;
			53756: outdata = 32'd11780;
			53757: outdata = 32'd11779;
			53758: outdata = 32'd11778;
			53759: outdata = 32'd11777;
			53760: outdata = 32'd11776;
			53761: outdata = 32'd11775;
			53762: outdata = 32'd11774;
			53763: outdata = 32'd11773;
			53764: outdata = 32'd11772;
			53765: outdata = 32'd11771;
			53766: outdata = 32'd11770;
			53767: outdata = 32'd11769;
			53768: outdata = 32'd11768;
			53769: outdata = 32'd11767;
			53770: outdata = 32'd11766;
			53771: outdata = 32'd11765;
			53772: outdata = 32'd11764;
			53773: outdata = 32'd11763;
			53774: outdata = 32'd11762;
			53775: outdata = 32'd11761;
			53776: outdata = 32'd11760;
			53777: outdata = 32'd11759;
			53778: outdata = 32'd11758;
			53779: outdata = 32'd11757;
			53780: outdata = 32'd11756;
			53781: outdata = 32'd11755;
			53782: outdata = 32'd11754;
			53783: outdata = 32'd11753;
			53784: outdata = 32'd11752;
			53785: outdata = 32'd11751;
			53786: outdata = 32'd11750;
			53787: outdata = 32'd11749;
			53788: outdata = 32'd11748;
			53789: outdata = 32'd11747;
			53790: outdata = 32'd11746;
			53791: outdata = 32'd11745;
			53792: outdata = 32'd11744;
			53793: outdata = 32'd11743;
			53794: outdata = 32'd11742;
			53795: outdata = 32'd11741;
			53796: outdata = 32'd11740;
			53797: outdata = 32'd11739;
			53798: outdata = 32'd11738;
			53799: outdata = 32'd11737;
			53800: outdata = 32'd11736;
			53801: outdata = 32'd11735;
			53802: outdata = 32'd11734;
			53803: outdata = 32'd11733;
			53804: outdata = 32'd11732;
			53805: outdata = 32'd11731;
			53806: outdata = 32'd11730;
			53807: outdata = 32'd11729;
			53808: outdata = 32'd11728;
			53809: outdata = 32'd11727;
			53810: outdata = 32'd11726;
			53811: outdata = 32'd11725;
			53812: outdata = 32'd11724;
			53813: outdata = 32'd11723;
			53814: outdata = 32'd11722;
			53815: outdata = 32'd11721;
			53816: outdata = 32'd11720;
			53817: outdata = 32'd11719;
			53818: outdata = 32'd11718;
			53819: outdata = 32'd11717;
			53820: outdata = 32'd11716;
			53821: outdata = 32'd11715;
			53822: outdata = 32'd11714;
			53823: outdata = 32'd11713;
			53824: outdata = 32'd11712;
			53825: outdata = 32'd11711;
			53826: outdata = 32'd11710;
			53827: outdata = 32'd11709;
			53828: outdata = 32'd11708;
			53829: outdata = 32'd11707;
			53830: outdata = 32'd11706;
			53831: outdata = 32'd11705;
			53832: outdata = 32'd11704;
			53833: outdata = 32'd11703;
			53834: outdata = 32'd11702;
			53835: outdata = 32'd11701;
			53836: outdata = 32'd11700;
			53837: outdata = 32'd11699;
			53838: outdata = 32'd11698;
			53839: outdata = 32'd11697;
			53840: outdata = 32'd11696;
			53841: outdata = 32'd11695;
			53842: outdata = 32'd11694;
			53843: outdata = 32'd11693;
			53844: outdata = 32'd11692;
			53845: outdata = 32'd11691;
			53846: outdata = 32'd11690;
			53847: outdata = 32'd11689;
			53848: outdata = 32'd11688;
			53849: outdata = 32'd11687;
			53850: outdata = 32'd11686;
			53851: outdata = 32'd11685;
			53852: outdata = 32'd11684;
			53853: outdata = 32'd11683;
			53854: outdata = 32'd11682;
			53855: outdata = 32'd11681;
			53856: outdata = 32'd11680;
			53857: outdata = 32'd11679;
			53858: outdata = 32'd11678;
			53859: outdata = 32'd11677;
			53860: outdata = 32'd11676;
			53861: outdata = 32'd11675;
			53862: outdata = 32'd11674;
			53863: outdata = 32'd11673;
			53864: outdata = 32'd11672;
			53865: outdata = 32'd11671;
			53866: outdata = 32'd11670;
			53867: outdata = 32'd11669;
			53868: outdata = 32'd11668;
			53869: outdata = 32'd11667;
			53870: outdata = 32'd11666;
			53871: outdata = 32'd11665;
			53872: outdata = 32'd11664;
			53873: outdata = 32'd11663;
			53874: outdata = 32'd11662;
			53875: outdata = 32'd11661;
			53876: outdata = 32'd11660;
			53877: outdata = 32'd11659;
			53878: outdata = 32'd11658;
			53879: outdata = 32'd11657;
			53880: outdata = 32'd11656;
			53881: outdata = 32'd11655;
			53882: outdata = 32'd11654;
			53883: outdata = 32'd11653;
			53884: outdata = 32'd11652;
			53885: outdata = 32'd11651;
			53886: outdata = 32'd11650;
			53887: outdata = 32'd11649;
			53888: outdata = 32'd11648;
			53889: outdata = 32'd11647;
			53890: outdata = 32'd11646;
			53891: outdata = 32'd11645;
			53892: outdata = 32'd11644;
			53893: outdata = 32'd11643;
			53894: outdata = 32'd11642;
			53895: outdata = 32'd11641;
			53896: outdata = 32'd11640;
			53897: outdata = 32'd11639;
			53898: outdata = 32'd11638;
			53899: outdata = 32'd11637;
			53900: outdata = 32'd11636;
			53901: outdata = 32'd11635;
			53902: outdata = 32'd11634;
			53903: outdata = 32'd11633;
			53904: outdata = 32'd11632;
			53905: outdata = 32'd11631;
			53906: outdata = 32'd11630;
			53907: outdata = 32'd11629;
			53908: outdata = 32'd11628;
			53909: outdata = 32'd11627;
			53910: outdata = 32'd11626;
			53911: outdata = 32'd11625;
			53912: outdata = 32'd11624;
			53913: outdata = 32'd11623;
			53914: outdata = 32'd11622;
			53915: outdata = 32'd11621;
			53916: outdata = 32'd11620;
			53917: outdata = 32'd11619;
			53918: outdata = 32'd11618;
			53919: outdata = 32'd11617;
			53920: outdata = 32'd11616;
			53921: outdata = 32'd11615;
			53922: outdata = 32'd11614;
			53923: outdata = 32'd11613;
			53924: outdata = 32'd11612;
			53925: outdata = 32'd11611;
			53926: outdata = 32'd11610;
			53927: outdata = 32'd11609;
			53928: outdata = 32'd11608;
			53929: outdata = 32'd11607;
			53930: outdata = 32'd11606;
			53931: outdata = 32'd11605;
			53932: outdata = 32'd11604;
			53933: outdata = 32'd11603;
			53934: outdata = 32'd11602;
			53935: outdata = 32'd11601;
			53936: outdata = 32'd11600;
			53937: outdata = 32'd11599;
			53938: outdata = 32'd11598;
			53939: outdata = 32'd11597;
			53940: outdata = 32'd11596;
			53941: outdata = 32'd11595;
			53942: outdata = 32'd11594;
			53943: outdata = 32'd11593;
			53944: outdata = 32'd11592;
			53945: outdata = 32'd11591;
			53946: outdata = 32'd11590;
			53947: outdata = 32'd11589;
			53948: outdata = 32'd11588;
			53949: outdata = 32'd11587;
			53950: outdata = 32'd11586;
			53951: outdata = 32'd11585;
			53952: outdata = 32'd11584;
			53953: outdata = 32'd11583;
			53954: outdata = 32'd11582;
			53955: outdata = 32'd11581;
			53956: outdata = 32'd11580;
			53957: outdata = 32'd11579;
			53958: outdata = 32'd11578;
			53959: outdata = 32'd11577;
			53960: outdata = 32'd11576;
			53961: outdata = 32'd11575;
			53962: outdata = 32'd11574;
			53963: outdata = 32'd11573;
			53964: outdata = 32'd11572;
			53965: outdata = 32'd11571;
			53966: outdata = 32'd11570;
			53967: outdata = 32'd11569;
			53968: outdata = 32'd11568;
			53969: outdata = 32'd11567;
			53970: outdata = 32'd11566;
			53971: outdata = 32'd11565;
			53972: outdata = 32'd11564;
			53973: outdata = 32'd11563;
			53974: outdata = 32'd11562;
			53975: outdata = 32'd11561;
			53976: outdata = 32'd11560;
			53977: outdata = 32'd11559;
			53978: outdata = 32'd11558;
			53979: outdata = 32'd11557;
			53980: outdata = 32'd11556;
			53981: outdata = 32'd11555;
			53982: outdata = 32'd11554;
			53983: outdata = 32'd11553;
			53984: outdata = 32'd11552;
			53985: outdata = 32'd11551;
			53986: outdata = 32'd11550;
			53987: outdata = 32'd11549;
			53988: outdata = 32'd11548;
			53989: outdata = 32'd11547;
			53990: outdata = 32'd11546;
			53991: outdata = 32'd11545;
			53992: outdata = 32'd11544;
			53993: outdata = 32'd11543;
			53994: outdata = 32'd11542;
			53995: outdata = 32'd11541;
			53996: outdata = 32'd11540;
			53997: outdata = 32'd11539;
			53998: outdata = 32'd11538;
			53999: outdata = 32'd11537;
			54000: outdata = 32'd11536;
			54001: outdata = 32'd11535;
			54002: outdata = 32'd11534;
			54003: outdata = 32'd11533;
			54004: outdata = 32'd11532;
			54005: outdata = 32'd11531;
			54006: outdata = 32'd11530;
			54007: outdata = 32'd11529;
			54008: outdata = 32'd11528;
			54009: outdata = 32'd11527;
			54010: outdata = 32'd11526;
			54011: outdata = 32'd11525;
			54012: outdata = 32'd11524;
			54013: outdata = 32'd11523;
			54014: outdata = 32'd11522;
			54015: outdata = 32'd11521;
			54016: outdata = 32'd11520;
			54017: outdata = 32'd11519;
			54018: outdata = 32'd11518;
			54019: outdata = 32'd11517;
			54020: outdata = 32'd11516;
			54021: outdata = 32'd11515;
			54022: outdata = 32'd11514;
			54023: outdata = 32'd11513;
			54024: outdata = 32'd11512;
			54025: outdata = 32'd11511;
			54026: outdata = 32'd11510;
			54027: outdata = 32'd11509;
			54028: outdata = 32'd11508;
			54029: outdata = 32'd11507;
			54030: outdata = 32'd11506;
			54031: outdata = 32'd11505;
			54032: outdata = 32'd11504;
			54033: outdata = 32'd11503;
			54034: outdata = 32'd11502;
			54035: outdata = 32'd11501;
			54036: outdata = 32'd11500;
			54037: outdata = 32'd11499;
			54038: outdata = 32'd11498;
			54039: outdata = 32'd11497;
			54040: outdata = 32'd11496;
			54041: outdata = 32'd11495;
			54042: outdata = 32'd11494;
			54043: outdata = 32'd11493;
			54044: outdata = 32'd11492;
			54045: outdata = 32'd11491;
			54046: outdata = 32'd11490;
			54047: outdata = 32'd11489;
			54048: outdata = 32'd11488;
			54049: outdata = 32'd11487;
			54050: outdata = 32'd11486;
			54051: outdata = 32'd11485;
			54052: outdata = 32'd11484;
			54053: outdata = 32'd11483;
			54054: outdata = 32'd11482;
			54055: outdata = 32'd11481;
			54056: outdata = 32'd11480;
			54057: outdata = 32'd11479;
			54058: outdata = 32'd11478;
			54059: outdata = 32'd11477;
			54060: outdata = 32'd11476;
			54061: outdata = 32'd11475;
			54062: outdata = 32'd11474;
			54063: outdata = 32'd11473;
			54064: outdata = 32'd11472;
			54065: outdata = 32'd11471;
			54066: outdata = 32'd11470;
			54067: outdata = 32'd11469;
			54068: outdata = 32'd11468;
			54069: outdata = 32'd11467;
			54070: outdata = 32'd11466;
			54071: outdata = 32'd11465;
			54072: outdata = 32'd11464;
			54073: outdata = 32'd11463;
			54074: outdata = 32'd11462;
			54075: outdata = 32'd11461;
			54076: outdata = 32'd11460;
			54077: outdata = 32'd11459;
			54078: outdata = 32'd11458;
			54079: outdata = 32'd11457;
			54080: outdata = 32'd11456;
			54081: outdata = 32'd11455;
			54082: outdata = 32'd11454;
			54083: outdata = 32'd11453;
			54084: outdata = 32'd11452;
			54085: outdata = 32'd11451;
			54086: outdata = 32'd11450;
			54087: outdata = 32'd11449;
			54088: outdata = 32'd11448;
			54089: outdata = 32'd11447;
			54090: outdata = 32'd11446;
			54091: outdata = 32'd11445;
			54092: outdata = 32'd11444;
			54093: outdata = 32'd11443;
			54094: outdata = 32'd11442;
			54095: outdata = 32'd11441;
			54096: outdata = 32'd11440;
			54097: outdata = 32'd11439;
			54098: outdata = 32'd11438;
			54099: outdata = 32'd11437;
			54100: outdata = 32'd11436;
			54101: outdata = 32'd11435;
			54102: outdata = 32'd11434;
			54103: outdata = 32'd11433;
			54104: outdata = 32'd11432;
			54105: outdata = 32'd11431;
			54106: outdata = 32'd11430;
			54107: outdata = 32'd11429;
			54108: outdata = 32'd11428;
			54109: outdata = 32'd11427;
			54110: outdata = 32'd11426;
			54111: outdata = 32'd11425;
			54112: outdata = 32'd11424;
			54113: outdata = 32'd11423;
			54114: outdata = 32'd11422;
			54115: outdata = 32'd11421;
			54116: outdata = 32'd11420;
			54117: outdata = 32'd11419;
			54118: outdata = 32'd11418;
			54119: outdata = 32'd11417;
			54120: outdata = 32'd11416;
			54121: outdata = 32'd11415;
			54122: outdata = 32'd11414;
			54123: outdata = 32'd11413;
			54124: outdata = 32'd11412;
			54125: outdata = 32'd11411;
			54126: outdata = 32'd11410;
			54127: outdata = 32'd11409;
			54128: outdata = 32'd11408;
			54129: outdata = 32'd11407;
			54130: outdata = 32'd11406;
			54131: outdata = 32'd11405;
			54132: outdata = 32'd11404;
			54133: outdata = 32'd11403;
			54134: outdata = 32'd11402;
			54135: outdata = 32'd11401;
			54136: outdata = 32'd11400;
			54137: outdata = 32'd11399;
			54138: outdata = 32'd11398;
			54139: outdata = 32'd11397;
			54140: outdata = 32'd11396;
			54141: outdata = 32'd11395;
			54142: outdata = 32'd11394;
			54143: outdata = 32'd11393;
			54144: outdata = 32'd11392;
			54145: outdata = 32'd11391;
			54146: outdata = 32'd11390;
			54147: outdata = 32'd11389;
			54148: outdata = 32'd11388;
			54149: outdata = 32'd11387;
			54150: outdata = 32'd11386;
			54151: outdata = 32'd11385;
			54152: outdata = 32'd11384;
			54153: outdata = 32'd11383;
			54154: outdata = 32'd11382;
			54155: outdata = 32'd11381;
			54156: outdata = 32'd11380;
			54157: outdata = 32'd11379;
			54158: outdata = 32'd11378;
			54159: outdata = 32'd11377;
			54160: outdata = 32'd11376;
			54161: outdata = 32'd11375;
			54162: outdata = 32'd11374;
			54163: outdata = 32'd11373;
			54164: outdata = 32'd11372;
			54165: outdata = 32'd11371;
			54166: outdata = 32'd11370;
			54167: outdata = 32'd11369;
			54168: outdata = 32'd11368;
			54169: outdata = 32'd11367;
			54170: outdata = 32'd11366;
			54171: outdata = 32'd11365;
			54172: outdata = 32'd11364;
			54173: outdata = 32'd11363;
			54174: outdata = 32'd11362;
			54175: outdata = 32'd11361;
			54176: outdata = 32'd11360;
			54177: outdata = 32'd11359;
			54178: outdata = 32'd11358;
			54179: outdata = 32'd11357;
			54180: outdata = 32'd11356;
			54181: outdata = 32'd11355;
			54182: outdata = 32'd11354;
			54183: outdata = 32'd11353;
			54184: outdata = 32'd11352;
			54185: outdata = 32'd11351;
			54186: outdata = 32'd11350;
			54187: outdata = 32'd11349;
			54188: outdata = 32'd11348;
			54189: outdata = 32'd11347;
			54190: outdata = 32'd11346;
			54191: outdata = 32'd11345;
			54192: outdata = 32'd11344;
			54193: outdata = 32'd11343;
			54194: outdata = 32'd11342;
			54195: outdata = 32'd11341;
			54196: outdata = 32'd11340;
			54197: outdata = 32'd11339;
			54198: outdata = 32'd11338;
			54199: outdata = 32'd11337;
			54200: outdata = 32'd11336;
			54201: outdata = 32'd11335;
			54202: outdata = 32'd11334;
			54203: outdata = 32'd11333;
			54204: outdata = 32'd11332;
			54205: outdata = 32'd11331;
			54206: outdata = 32'd11330;
			54207: outdata = 32'd11329;
			54208: outdata = 32'd11328;
			54209: outdata = 32'd11327;
			54210: outdata = 32'd11326;
			54211: outdata = 32'd11325;
			54212: outdata = 32'd11324;
			54213: outdata = 32'd11323;
			54214: outdata = 32'd11322;
			54215: outdata = 32'd11321;
			54216: outdata = 32'd11320;
			54217: outdata = 32'd11319;
			54218: outdata = 32'd11318;
			54219: outdata = 32'd11317;
			54220: outdata = 32'd11316;
			54221: outdata = 32'd11315;
			54222: outdata = 32'd11314;
			54223: outdata = 32'd11313;
			54224: outdata = 32'd11312;
			54225: outdata = 32'd11311;
			54226: outdata = 32'd11310;
			54227: outdata = 32'd11309;
			54228: outdata = 32'd11308;
			54229: outdata = 32'd11307;
			54230: outdata = 32'd11306;
			54231: outdata = 32'd11305;
			54232: outdata = 32'd11304;
			54233: outdata = 32'd11303;
			54234: outdata = 32'd11302;
			54235: outdata = 32'd11301;
			54236: outdata = 32'd11300;
			54237: outdata = 32'd11299;
			54238: outdata = 32'd11298;
			54239: outdata = 32'd11297;
			54240: outdata = 32'd11296;
			54241: outdata = 32'd11295;
			54242: outdata = 32'd11294;
			54243: outdata = 32'd11293;
			54244: outdata = 32'd11292;
			54245: outdata = 32'd11291;
			54246: outdata = 32'd11290;
			54247: outdata = 32'd11289;
			54248: outdata = 32'd11288;
			54249: outdata = 32'd11287;
			54250: outdata = 32'd11286;
			54251: outdata = 32'd11285;
			54252: outdata = 32'd11284;
			54253: outdata = 32'd11283;
			54254: outdata = 32'd11282;
			54255: outdata = 32'd11281;
			54256: outdata = 32'd11280;
			54257: outdata = 32'd11279;
			54258: outdata = 32'd11278;
			54259: outdata = 32'd11277;
			54260: outdata = 32'd11276;
			54261: outdata = 32'd11275;
			54262: outdata = 32'd11274;
			54263: outdata = 32'd11273;
			54264: outdata = 32'd11272;
			54265: outdata = 32'd11271;
			54266: outdata = 32'd11270;
			54267: outdata = 32'd11269;
			54268: outdata = 32'd11268;
			54269: outdata = 32'd11267;
			54270: outdata = 32'd11266;
			54271: outdata = 32'd11265;
			54272: outdata = 32'd11264;
			54273: outdata = 32'd11263;
			54274: outdata = 32'd11262;
			54275: outdata = 32'd11261;
			54276: outdata = 32'd11260;
			54277: outdata = 32'd11259;
			54278: outdata = 32'd11258;
			54279: outdata = 32'd11257;
			54280: outdata = 32'd11256;
			54281: outdata = 32'd11255;
			54282: outdata = 32'd11254;
			54283: outdata = 32'd11253;
			54284: outdata = 32'd11252;
			54285: outdata = 32'd11251;
			54286: outdata = 32'd11250;
			54287: outdata = 32'd11249;
			54288: outdata = 32'd11248;
			54289: outdata = 32'd11247;
			54290: outdata = 32'd11246;
			54291: outdata = 32'd11245;
			54292: outdata = 32'd11244;
			54293: outdata = 32'd11243;
			54294: outdata = 32'd11242;
			54295: outdata = 32'd11241;
			54296: outdata = 32'd11240;
			54297: outdata = 32'd11239;
			54298: outdata = 32'd11238;
			54299: outdata = 32'd11237;
			54300: outdata = 32'd11236;
			54301: outdata = 32'd11235;
			54302: outdata = 32'd11234;
			54303: outdata = 32'd11233;
			54304: outdata = 32'd11232;
			54305: outdata = 32'd11231;
			54306: outdata = 32'd11230;
			54307: outdata = 32'd11229;
			54308: outdata = 32'd11228;
			54309: outdata = 32'd11227;
			54310: outdata = 32'd11226;
			54311: outdata = 32'd11225;
			54312: outdata = 32'd11224;
			54313: outdata = 32'd11223;
			54314: outdata = 32'd11222;
			54315: outdata = 32'd11221;
			54316: outdata = 32'd11220;
			54317: outdata = 32'd11219;
			54318: outdata = 32'd11218;
			54319: outdata = 32'd11217;
			54320: outdata = 32'd11216;
			54321: outdata = 32'd11215;
			54322: outdata = 32'd11214;
			54323: outdata = 32'd11213;
			54324: outdata = 32'd11212;
			54325: outdata = 32'd11211;
			54326: outdata = 32'd11210;
			54327: outdata = 32'd11209;
			54328: outdata = 32'd11208;
			54329: outdata = 32'd11207;
			54330: outdata = 32'd11206;
			54331: outdata = 32'd11205;
			54332: outdata = 32'd11204;
			54333: outdata = 32'd11203;
			54334: outdata = 32'd11202;
			54335: outdata = 32'd11201;
			54336: outdata = 32'd11200;
			54337: outdata = 32'd11199;
			54338: outdata = 32'd11198;
			54339: outdata = 32'd11197;
			54340: outdata = 32'd11196;
			54341: outdata = 32'd11195;
			54342: outdata = 32'd11194;
			54343: outdata = 32'd11193;
			54344: outdata = 32'd11192;
			54345: outdata = 32'd11191;
			54346: outdata = 32'd11190;
			54347: outdata = 32'd11189;
			54348: outdata = 32'd11188;
			54349: outdata = 32'd11187;
			54350: outdata = 32'd11186;
			54351: outdata = 32'd11185;
			54352: outdata = 32'd11184;
			54353: outdata = 32'd11183;
			54354: outdata = 32'd11182;
			54355: outdata = 32'd11181;
			54356: outdata = 32'd11180;
			54357: outdata = 32'd11179;
			54358: outdata = 32'd11178;
			54359: outdata = 32'd11177;
			54360: outdata = 32'd11176;
			54361: outdata = 32'd11175;
			54362: outdata = 32'd11174;
			54363: outdata = 32'd11173;
			54364: outdata = 32'd11172;
			54365: outdata = 32'd11171;
			54366: outdata = 32'd11170;
			54367: outdata = 32'd11169;
			54368: outdata = 32'd11168;
			54369: outdata = 32'd11167;
			54370: outdata = 32'd11166;
			54371: outdata = 32'd11165;
			54372: outdata = 32'd11164;
			54373: outdata = 32'd11163;
			54374: outdata = 32'd11162;
			54375: outdata = 32'd11161;
			54376: outdata = 32'd11160;
			54377: outdata = 32'd11159;
			54378: outdata = 32'd11158;
			54379: outdata = 32'd11157;
			54380: outdata = 32'd11156;
			54381: outdata = 32'd11155;
			54382: outdata = 32'd11154;
			54383: outdata = 32'd11153;
			54384: outdata = 32'd11152;
			54385: outdata = 32'd11151;
			54386: outdata = 32'd11150;
			54387: outdata = 32'd11149;
			54388: outdata = 32'd11148;
			54389: outdata = 32'd11147;
			54390: outdata = 32'd11146;
			54391: outdata = 32'd11145;
			54392: outdata = 32'd11144;
			54393: outdata = 32'd11143;
			54394: outdata = 32'd11142;
			54395: outdata = 32'd11141;
			54396: outdata = 32'd11140;
			54397: outdata = 32'd11139;
			54398: outdata = 32'd11138;
			54399: outdata = 32'd11137;
			54400: outdata = 32'd11136;
			54401: outdata = 32'd11135;
			54402: outdata = 32'd11134;
			54403: outdata = 32'd11133;
			54404: outdata = 32'd11132;
			54405: outdata = 32'd11131;
			54406: outdata = 32'd11130;
			54407: outdata = 32'd11129;
			54408: outdata = 32'd11128;
			54409: outdata = 32'd11127;
			54410: outdata = 32'd11126;
			54411: outdata = 32'd11125;
			54412: outdata = 32'd11124;
			54413: outdata = 32'd11123;
			54414: outdata = 32'd11122;
			54415: outdata = 32'd11121;
			54416: outdata = 32'd11120;
			54417: outdata = 32'd11119;
			54418: outdata = 32'd11118;
			54419: outdata = 32'd11117;
			54420: outdata = 32'd11116;
			54421: outdata = 32'd11115;
			54422: outdata = 32'd11114;
			54423: outdata = 32'd11113;
			54424: outdata = 32'd11112;
			54425: outdata = 32'd11111;
			54426: outdata = 32'd11110;
			54427: outdata = 32'd11109;
			54428: outdata = 32'd11108;
			54429: outdata = 32'd11107;
			54430: outdata = 32'd11106;
			54431: outdata = 32'd11105;
			54432: outdata = 32'd11104;
			54433: outdata = 32'd11103;
			54434: outdata = 32'd11102;
			54435: outdata = 32'd11101;
			54436: outdata = 32'd11100;
			54437: outdata = 32'd11099;
			54438: outdata = 32'd11098;
			54439: outdata = 32'd11097;
			54440: outdata = 32'd11096;
			54441: outdata = 32'd11095;
			54442: outdata = 32'd11094;
			54443: outdata = 32'd11093;
			54444: outdata = 32'd11092;
			54445: outdata = 32'd11091;
			54446: outdata = 32'd11090;
			54447: outdata = 32'd11089;
			54448: outdata = 32'd11088;
			54449: outdata = 32'd11087;
			54450: outdata = 32'd11086;
			54451: outdata = 32'd11085;
			54452: outdata = 32'd11084;
			54453: outdata = 32'd11083;
			54454: outdata = 32'd11082;
			54455: outdata = 32'd11081;
			54456: outdata = 32'd11080;
			54457: outdata = 32'd11079;
			54458: outdata = 32'd11078;
			54459: outdata = 32'd11077;
			54460: outdata = 32'd11076;
			54461: outdata = 32'd11075;
			54462: outdata = 32'd11074;
			54463: outdata = 32'd11073;
			54464: outdata = 32'd11072;
			54465: outdata = 32'd11071;
			54466: outdata = 32'd11070;
			54467: outdata = 32'd11069;
			54468: outdata = 32'd11068;
			54469: outdata = 32'd11067;
			54470: outdata = 32'd11066;
			54471: outdata = 32'd11065;
			54472: outdata = 32'd11064;
			54473: outdata = 32'd11063;
			54474: outdata = 32'd11062;
			54475: outdata = 32'd11061;
			54476: outdata = 32'd11060;
			54477: outdata = 32'd11059;
			54478: outdata = 32'd11058;
			54479: outdata = 32'd11057;
			54480: outdata = 32'd11056;
			54481: outdata = 32'd11055;
			54482: outdata = 32'd11054;
			54483: outdata = 32'd11053;
			54484: outdata = 32'd11052;
			54485: outdata = 32'd11051;
			54486: outdata = 32'd11050;
			54487: outdata = 32'd11049;
			54488: outdata = 32'd11048;
			54489: outdata = 32'd11047;
			54490: outdata = 32'd11046;
			54491: outdata = 32'd11045;
			54492: outdata = 32'd11044;
			54493: outdata = 32'd11043;
			54494: outdata = 32'd11042;
			54495: outdata = 32'd11041;
			54496: outdata = 32'd11040;
			54497: outdata = 32'd11039;
			54498: outdata = 32'd11038;
			54499: outdata = 32'd11037;
			54500: outdata = 32'd11036;
			54501: outdata = 32'd11035;
			54502: outdata = 32'd11034;
			54503: outdata = 32'd11033;
			54504: outdata = 32'd11032;
			54505: outdata = 32'd11031;
			54506: outdata = 32'd11030;
			54507: outdata = 32'd11029;
			54508: outdata = 32'd11028;
			54509: outdata = 32'd11027;
			54510: outdata = 32'd11026;
			54511: outdata = 32'd11025;
			54512: outdata = 32'd11024;
			54513: outdata = 32'd11023;
			54514: outdata = 32'd11022;
			54515: outdata = 32'd11021;
			54516: outdata = 32'd11020;
			54517: outdata = 32'd11019;
			54518: outdata = 32'd11018;
			54519: outdata = 32'd11017;
			54520: outdata = 32'd11016;
			54521: outdata = 32'd11015;
			54522: outdata = 32'd11014;
			54523: outdata = 32'd11013;
			54524: outdata = 32'd11012;
			54525: outdata = 32'd11011;
			54526: outdata = 32'd11010;
			54527: outdata = 32'd11009;
			54528: outdata = 32'd11008;
			54529: outdata = 32'd11007;
			54530: outdata = 32'd11006;
			54531: outdata = 32'd11005;
			54532: outdata = 32'd11004;
			54533: outdata = 32'd11003;
			54534: outdata = 32'd11002;
			54535: outdata = 32'd11001;
			54536: outdata = 32'd11000;
			54537: outdata = 32'd10999;
			54538: outdata = 32'd10998;
			54539: outdata = 32'd10997;
			54540: outdata = 32'd10996;
			54541: outdata = 32'd10995;
			54542: outdata = 32'd10994;
			54543: outdata = 32'd10993;
			54544: outdata = 32'd10992;
			54545: outdata = 32'd10991;
			54546: outdata = 32'd10990;
			54547: outdata = 32'd10989;
			54548: outdata = 32'd10988;
			54549: outdata = 32'd10987;
			54550: outdata = 32'd10986;
			54551: outdata = 32'd10985;
			54552: outdata = 32'd10984;
			54553: outdata = 32'd10983;
			54554: outdata = 32'd10982;
			54555: outdata = 32'd10981;
			54556: outdata = 32'd10980;
			54557: outdata = 32'd10979;
			54558: outdata = 32'd10978;
			54559: outdata = 32'd10977;
			54560: outdata = 32'd10976;
			54561: outdata = 32'd10975;
			54562: outdata = 32'd10974;
			54563: outdata = 32'd10973;
			54564: outdata = 32'd10972;
			54565: outdata = 32'd10971;
			54566: outdata = 32'd10970;
			54567: outdata = 32'd10969;
			54568: outdata = 32'd10968;
			54569: outdata = 32'd10967;
			54570: outdata = 32'd10966;
			54571: outdata = 32'd10965;
			54572: outdata = 32'd10964;
			54573: outdata = 32'd10963;
			54574: outdata = 32'd10962;
			54575: outdata = 32'd10961;
			54576: outdata = 32'd10960;
			54577: outdata = 32'd10959;
			54578: outdata = 32'd10958;
			54579: outdata = 32'd10957;
			54580: outdata = 32'd10956;
			54581: outdata = 32'd10955;
			54582: outdata = 32'd10954;
			54583: outdata = 32'd10953;
			54584: outdata = 32'd10952;
			54585: outdata = 32'd10951;
			54586: outdata = 32'd10950;
			54587: outdata = 32'd10949;
			54588: outdata = 32'd10948;
			54589: outdata = 32'd10947;
			54590: outdata = 32'd10946;
			54591: outdata = 32'd10945;
			54592: outdata = 32'd10944;
			54593: outdata = 32'd10943;
			54594: outdata = 32'd10942;
			54595: outdata = 32'd10941;
			54596: outdata = 32'd10940;
			54597: outdata = 32'd10939;
			54598: outdata = 32'd10938;
			54599: outdata = 32'd10937;
			54600: outdata = 32'd10936;
			54601: outdata = 32'd10935;
			54602: outdata = 32'd10934;
			54603: outdata = 32'd10933;
			54604: outdata = 32'd10932;
			54605: outdata = 32'd10931;
			54606: outdata = 32'd10930;
			54607: outdata = 32'd10929;
			54608: outdata = 32'd10928;
			54609: outdata = 32'd10927;
			54610: outdata = 32'd10926;
			54611: outdata = 32'd10925;
			54612: outdata = 32'd10924;
			54613: outdata = 32'd10923;
			54614: outdata = 32'd10922;
			54615: outdata = 32'd10921;
			54616: outdata = 32'd10920;
			54617: outdata = 32'd10919;
			54618: outdata = 32'd10918;
			54619: outdata = 32'd10917;
			54620: outdata = 32'd10916;
			54621: outdata = 32'd10915;
			54622: outdata = 32'd10914;
			54623: outdata = 32'd10913;
			54624: outdata = 32'd10912;
			54625: outdata = 32'd10911;
			54626: outdata = 32'd10910;
			54627: outdata = 32'd10909;
			54628: outdata = 32'd10908;
			54629: outdata = 32'd10907;
			54630: outdata = 32'd10906;
			54631: outdata = 32'd10905;
			54632: outdata = 32'd10904;
			54633: outdata = 32'd10903;
			54634: outdata = 32'd10902;
			54635: outdata = 32'd10901;
			54636: outdata = 32'd10900;
			54637: outdata = 32'd10899;
			54638: outdata = 32'd10898;
			54639: outdata = 32'd10897;
			54640: outdata = 32'd10896;
			54641: outdata = 32'd10895;
			54642: outdata = 32'd10894;
			54643: outdata = 32'd10893;
			54644: outdata = 32'd10892;
			54645: outdata = 32'd10891;
			54646: outdata = 32'd10890;
			54647: outdata = 32'd10889;
			54648: outdata = 32'd10888;
			54649: outdata = 32'd10887;
			54650: outdata = 32'd10886;
			54651: outdata = 32'd10885;
			54652: outdata = 32'd10884;
			54653: outdata = 32'd10883;
			54654: outdata = 32'd10882;
			54655: outdata = 32'd10881;
			54656: outdata = 32'd10880;
			54657: outdata = 32'd10879;
			54658: outdata = 32'd10878;
			54659: outdata = 32'd10877;
			54660: outdata = 32'd10876;
			54661: outdata = 32'd10875;
			54662: outdata = 32'd10874;
			54663: outdata = 32'd10873;
			54664: outdata = 32'd10872;
			54665: outdata = 32'd10871;
			54666: outdata = 32'd10870;
			54667: outdata = 32'd10869;
			54668: outdata = 32'd10868;
			54669: outdata = 32'd10867;
			54670: outdata = 32'd10866;
			54671: outdata = 32'd10865;
			54672: outdata = 32'd10864;
			54673: outdata = 32'd10863;
			54674: outdata = 32'd10862;
			54675: outdata = 32'd10861;
			54676: outdata = 32'd10860;
			54677: outdata = 32'd10859;
			54678: outdata = 32'd10858;
			54679: outdata = 32'd10857;
			54680: outdata = 32'd10856;
			54681: outdata = 32'd10855;
			54682: outdata = 32'd10854;
			54683: outdata = 32'd10853;
			54684: outdata = 32'd10852;
			54685: outdata = 32'd10851;
			54686: outdata = 32'd10850;
			54687: outdata = 32'd10849;
			54688: outdata = 32'd10848;
			54689: outdata = 32'd10847;
			54690: outdata = 32'd10846;
			54691: outdata = 32'd10845;
			54692: outdata = 32'd10844;
			54693: outdata = 32'd10843;
			54694: outdata = 32'd10842;
			54695: outdata = 32'd10841;
			54696: outdata = 32'd10840;
			54697: outdata = 32'd10839;
			54698: outdata = 32'd10838;
			54699: outdata = 32'd10837;
			54700: outdata = 32'd10836;
			54701: outdata = 32'd10835;
			54702: outdata = 32'd10834;
			54703: outdata = 32'd10833;
			54704: outdata = 32'd10832;
			54705: outdata = 32'd10831;
			54706: outdata = 32'd10830;
			54707: outdata = 32'd10829;
			54708: outdata = 32'd10828;
			54709: outdata = 32'd10827;
			54710: outdata = 32'd10826;
			54711: outdata = 32'd10825;
			54712: outdata = 32'd10824;
			54713: outdata = 32'd10823;
			54714: outdata = 32'd10822;
			54715: outdata = 32'd10821;
			54716: outdata = 32'd10820;
			54717: outdata = 32'd10819;
			54718: outdata = 32'd10818;
			54719: outdata = 32'd10817;
			54720: outdata = 32'd10816;
			54721: outdata = 32'd10815;
			54722: outdata = 32'd10814;
			54723: outdata = 32'd10813;
			54724: outdata = 32'd10812;
			54725: outdata = 32'd10811;
			54726: outdata = 32'd10810;
			54727: outdata = 32'd10809;
			54728: outdata = 32'd10808;
			54729: outdata = 32'd10807;
			54730: outdata = 32'd10806;
			54731: outdata = 32'd10805;
			54732: outdata = 32'd10804;
			54733: outdata = 32'd10803;
			54734: outdata = 32'd10802;
			54735: outdata = 32'd10801;
			54736: outdata = 32'd10800;
			54737: outdata = 32'd10799;
			54738: outdata = 32'd10798;
			54739: outdata = 32'd10797;
			54740: outdata = 32'd10796;
			54741: outdata = 32'd10795;
			54742: outdata = 32'd10794;
			54743: outdata = 32'd10793;
			54744: outdata = 32'd10792;
			54745: outdata = 32'd10791;
			54746: outdata = 32'd10790;
			54747: outdata = 32'd10789;
			54748: outdata = 32'd10788;
			54749: outdata = 32'd10787;
			54750: outdata = 32'd10786;
			54751: outdata = 32'd10785;
			54752: outdata = 32'd10784;
			54753: outdata = 32'd10783;
			54754: outdata = 32'd10782;
			54755: outdata = 32'd10781;
			54756: outdata = 32'd10780;
			54757: outdata = 32'd10779;
			54758: outdata = 32'd10778;
			54759: outdata = 32'd10777;
			54760: outdata = 32'd10776;
			54761: outdata = 32'd10775;
			54762: outdata = 32'd10774;
			54763: outdata = 32'd10773;
			54764: outdata = 32'd10772;
			54765: outdata = 32'd10771;
			54766: outdata = 32'd10770;
			54767: outdata = 32'd10769;
			54768: outdata = 32'd10768;
			54769: outdata = 32'd10767;
			54770: outdata = 32'd10766;
			54771: outdata = 32'd10765;
			54772: outdata = 32'd10764;
			54773: outdata = 32'd10763;
			54774: outdata = 32'd10762;
			54775: outdata = 32'd10761;
			54776: outdata = 32'd10760;
			54777: outdata = 32'd10759;
			54778: outdata = 32'd10758;
			54779: outdata = 32'd10757;
			54780: outdata = 32'd10756;
			54781: outdata = 32'd10755;
			54782: outdata = 32'd10754;
			54783: outdata = 32'd10753;
			54784: outdata = 32'd10752;
			54785: outdata = 32'd10751;
			54786: outdata = 32'd10750;
			54787: outdata = 32'd10749;
			54788: outdata = 32'd10748;
			54789: outdata = 32'd10747;
			54790: outdata = 32'd10746;
			54791: outdata = 32'd10745;
			54792: outdata = 32'd10744;
			54793: outdata = 32'd10743;
			54794: outdata = 32'd10742;
			54795: outdata = 32'd10741;
			54796: outdata = 32'd10740;
			54797: outdata = 32'd10739;
			54798: outdata = 32'd10738;
			54799: outdata = 32'd10737;
			54800: outdata = 32'd10736;
			54801: outdata = 32'd10735;
			54802: outdata = 32'd10734;
			54803: outdata = 32'd10733;
			54804: outdata = 32'd10732;
			54805: outdata = 32'd10731;
			54806: outdata = 32'd10730;
			54807: outdata = 32'd10729;
			54808: outdata = 32'd10728;
			54809: outdata = 32'd10727;
			54810: outdata = 32'd10726;
			54811: outdata = 32'd10725;
			54812: outdata = 32'd10724;
			54813: outdata = 32'd10723;
			54814: outdata = 32'd10722;
			54815: outdata = 32'd10721;
			54816: outdata = 32'd10720;
			54817: outdata = 32'd10719;
			54818: outdata = 32'd10718;
			54819: outdata = 32'd10717;
			54820: outdata = 32'd10716;
			54821: outdata = 32'd10715;
			54822: outdata = 32'd10714;
			54823: outdata = 32'd10713;
			54824: outdata = 32'd10712;
			54825: outdata = 32'd10711;
			54826: outdata = 32'd10710;
			54827: outdata = 32'd10709;
			54828: outdata = 32'd10708;
			54829: outdata = 32'd10707;
			54830: outdata = 32'd10706;
			54831: outdata = 32'd10705;
			54832: outdata = 32'd10704;
			54833: outdata = 32'd10703;
			54834: outdata = 32'd10702;
			54835: outdata = 32'd10701;
			54836: outdata = 32'd10700;
			54837: outdata = 32'd10699;
			54838: outdata = 32'd10698;
			54839: outdata = 32'd10697;
			54840: outdata = 32'd10696;
			54841: outdata = 32'd10695;
			54842: outdata = 32'd10694;
			54843: outdata = 32'd10693;
			54844: outdata = 32'd10692;
			54845: outdata = 32'd10691;
			54846: outdata = 32'd10690;
			54847: outdata = 32'd10689;
			54848: outdata = 32'd10688;
			54849: outdata = 32'd10687;
			54850: outdata = 32'd10686;
			54851: outdata = 32'd10685;
			54852: outdata = 32'd10684;
			54853: outdata = 32'd10683;
			54854: outdata = 32'd10682;
			54855: outdata = 32'd10681;
			54856: outdata = 32'd10680;
			54857: outdata = 32'd10679;
			54858: outdata = 32'd10678;
			54859: outdata = 32'd10677;
			54860: outdata = 32'd10676;
			54861: outdata = 32'd10675;
			54862: outdata = 32'd10674;
			54863: outdata = 32'd10673;
			54864: outdata = 32'd10672;
			54865: outdata = 32'd10671;
			54866: outdata = 32'd10670;
			54867: outdata = 32'd10669;
			54868: outdata = 32'd10668;
			54869: outdata = 32'd10667;
			54870: outdata = 32'd10666;
			54871: outdata = 32'd10665;
			54872: outdata = 32'd10664;
			54873: outdata = 32'd10663;
			54874: outdata = 32'd10662;
			54875: outdata = 32'd10661;
			54876: outdata = 32'd10660;
			54877: outdata = 32'd10659;
			54878: outdata = 32'd10658;
			54879: outdata = 32'd10657;
			54880: outdata = 32'd10656;
			54881: outdata = 32'd10655;
			54882: outdata = 32'd10654;
			54883: outdata = 32'd10653;
			54884: outdata = 32'd10652;
			54885: outdata = 32'd10651;
			54886: outdata = 32'd10650;
			54887: outdata = 32'd10649;
			54888: outdata = 32'd10648;
			54889: outdata = 32'd10647;
			54890: outdata = 32'd10646;
			54891: outdata = 32'd10645;
			54892: outdata = 32'd10644;
			54893: outdata = 32'd10643;
			54894: outdata = 32'd10642;
			54895: outdata = 32'd10641;
			54896: outdata = 32'd10640;
			54897: outdata = 32'd10639;
			54898: outdata = 32'd10638;
			54899: outdata = 32'd10637;
			54900: outdata = 32'd10636;
			54901: outdata = 32'd10635;
			54902: outdata = 32'd10634;
			54903: outdata = 32'd10633;
			54904: outdata = 32'd10632;
			54905: outdata = 32'd10631;
			54906: outdata = 32'd10630;
			54907: outdata = 32'd10629;
			54908: outdata = 32'd10628;
			54909: outdata = 32'd10627;
			54910: outdata = 32'd10626;
			54911: outdata = 32'd10625;
			54912: outdata = 32'd10624;
			54913: outdata = 32'd10623;
			54914: outdata = 32'd10622;
			54915: outdata = 32'd10621;
			54916: outdata = 32'd10620;
			54917: outdata = 32'd10619;
			54918: outdata = 32'd10618;
			54919: outdata = 32'd10617;
			54920: outdata = 32'd10616;
			54921: outdata = 32'd10615;
			54922: outdata = 32'd10614;
			54923: outdata = 32'd10613;
			54924: outdata = 32'd10612;
			54925: outdata = 32'd10611;
			54926: outdata = 32'd10610;
			54927: outdata = 32'd10609;
			54928: outdata = 32'd10608;
			54929: outdata = 32'd10607;
			54930: outdata = 32'd10606;
			54931: outdata = 32'd10605;
			54932: outdata = 32'd10604;
			54933: outdata = 32'd10603;
			54934: outdata = 32'd10602;
			54935: outdata = 32'd10601;
			54936: outdata = 32'd10600;
			54937: outdata = 32'd10599;
			54938: outdata = 32'd10598;
			54939: outdata = 32'd10597;
			54940: outdata = 32'd10596;
			54941: outdata = 32'd10595;
			54942: outdata = 32'd10594;
			54943: outdata = 32'd10593;
			54944: outdata = 32'd10592;
			54945: outdata = 32'd10591;
			54946: outdata = 32'd10590;
			54947: outdata = 32'd10589;
			54948: outdata = 32'd10588;
			54949: outdata = 32'd10587;
			54950: outdata = 32'd10586;
			54951: outdata = 32'd10585;
			54952: outdata = 32'd10584;
			54953: outdata = 32'd10583;
			54954: outdata = 32'd10582;
			54955: outdata = 32'd10581;
			54956: outdata = 32'd10580;
			54957: outdata = 32'd10579;
			54958: outdata = 32'd10578;
			54959: outdata = 32'd10577;
			54960: outdata = 32'd10576;
			54961: outdata = 32'd10575;
			54962: outdata = 32'd10574;
			54963: outdata = 32'd10573;
			54964: outdata = 32'd10572;
			54965: outdata = 32'd10571;
			54966: outdata = 32'd10570;
			54967: outdata = 32'd10569;
			54968: outdata = 32'd10568;
			54969: outdata = 32'd10567;
			54970: outdata = 32'd10566;
			54971: outdata = 32'd10565;
			54972: outdata = 32'd10564;
			54973: outdata = 32'd10563;
			54974: outdata = 32'd10562;
			54975: outdata = 32'd10561;
			54976: outdata = 32'd10560;
			54977: outdata = 32'd10559;
			54978: outdata = 32'd10558;
			54979: outdata = 32'd10557;
			54980: outdata = 32'd10556;
			54981: outdata = 32'd10555;
			54982: outdata = 32'd10554;
			54983: outdata = 32'd10553;
			54984: outdata = 32'd10552;
			54985: outdata = 32'd10551;
			54986: outdata = 32'd10550;
			54987: outdata = 32'd10549;
			54988: outdata = 32'd10548;
			54989: outdata = 32'd10547;
			54990: outdata = 32'd10546;
			54991: outdata = 32'd10545;
			54992: outdata = 32'd10544;
			54993: outdata = 32'd10543;
			54994: outdata = 32'd10542;
			54995: outdata = 32'd10541;
			54996: outdata = 32'd10540;
			54997: outdata = 32'd10539;
			54998: outdata = 32'd10538;
			54999: outdata = 32'd10537;
			55000: outdata = 32'd10536;
			55001: outdata = 32'd10535;
			55002: outdata = 32'd10534;
			55003: outdata = 32'd10533;
			55004: outdata = 32'd10532;
			55005: outdata = 32'd10531;
			55006: outdata = 32'd10530;
			55007: outdata = 32'd10529;
			55008: outdata = 32'd10528;
			55009: outdata = 32'd10527;
			55010: outdata = 32'd10526;
			55011: outdata = 32'd10525;
			55012: outdata = 32'd10524;
			55013: outdata = 32'd10523;
			55014: outdata = 32'd10522;
			55015: outdata = 32'd10521;
			55016: outdata = 32'd10520;
			55017: outdata = 32'd10519;
			55018: outdata = 32'd10518;
			55019: outdata = 32'd10517;
			55020: outdata = 32'd10516;
			55021: outdata = 32'd10515;
			55022: outdata = 32'd10514;
			55023: outdata = 32'd10513;
			55024: outdata = 32'd10512;
			55025: outdata = 32'd10511;
			55026: outdata = 32'd10510;
			55027: outdata = 32'd10509;
			55028: outdata = 32'd10508;
			55029: outdata = 32'd10507;
			55030: outdata = 32'd10506;
			55031: outdata = 32'd10505;
			55032: outdata = 32'd10504;
			55033: outdata = 32'd10503;
			55034: outdata = 32'd10502;
			55035: outdata = 32'd10501;
			55036: outdata = 32'd10500;
			55037: outdata = 32'd10499;
			55038: outdata = 32'd10498;
			55039: outdata = 32'd10497;
			55040: outdata = 32'd10496;
			55041: outdata = 32'd10495;
			55042: outdata = 32'd10494;
			55043: outdata = 32'd10493;
			55044: outdata = 32'd10492;
			55045: outdata = 32'd10491;
			55046: outdata = 32'd10490;
			55047: outdata = 32'd10489;
			55048: outdata = 32'd10488;
			55049: outdata = 32'd10487;
			55050: outdata = 32'd10486;
			55051: outdata = 32'd10485;
			55052: outdata = 32'd10484;
			55053: outdata = 32'd10483;
			55054: outdata = 32'd10482;
			55055: outdata = 32'd10481;
			55056: outdata = 32'd10480;
			55057: outdata = 32'd10479;
			55058: outdata = 32'd10478;
			55059: outdata = 32'd10477;
			55060: outdata = 32'd10476;
			55061: outdata = 32'd10475;
			55062: outdata = 32'd10474;
			55063: outdata = 32'd10473;
			55064: outdata = 32'd10472;
			55065: outdata = 32'd10471;
			55066: outdata = 32'd10470;
			55067: outdata = 32'd10469;
			55068: outdata = 32'd10468;
			55069: outdata = 32'd10467;
			55070: outdata = 32'd10466;
			55071: outdata = 32'd10465;
			55072: outdata = 32'd10464;
			55073: outdata = 32'd10463;
			55074: outdata = 32'd10462;
			55075: outdata = 32'd10461;
			55076: outdata = 32'd10460;
			55077: outdata = 32'd10459;
			55078: outdata = 32'd10458;
			55079: outdata = 32'd10457;
			55080: outdata = 32'd10456;
			55081: outdata = 32'd10455;
			55082: outdata = 32'd10454;
			55083: outdata = 32'd10453;
			55084: outdata = 32'd10452;
			55085: outdata = 32'd10451;
			55086: outdata = 32'd10450;
			55087: outdata = 32'd10449;
			55088: outdata = 32'd10448;
			55089: outdata = 32'd10447;
			55090: outdata = 32'd10446;
			55091: outdata = 32'd10445;
			55092: outdata = 32'd10444;
			55093: outdata = 32'd10443;
			55094: outdata = 32'd10442;
			55095: outdata = 32'd10441;
			55096: outdata = 32'd10440;
			55097: outdata = 32'd10439;
			55098: outdata = 32'd10438;
			55099: outdata = 32'd10437;
			55100: outdata = 32'd10436;
			55101: outdata = 32'd10435;
			55102: outdata = 32'd10434;
			55103: outdata = 32'd10433;
			55104: outdata = 32'd10432;
			55105: outdata = 32'd10431;
			55106: outdata = 32'd10430;
			55107: outdata = 32'd10429;
			55108: outdata = 32'd10428;
			55109: outdata = 32'd10427;
			55110: outdata = 32'd10426;
			55111: outdata = 32'd10425;
			55112: outdata = 32'd10424;
			55113: outdata = 32'd10423;
			55114: outdata = 32'd10422;
			55115: outdata = 32'd10421;
			55116: outdata = 32'd10420;
			55117: outdata = 32'd10419;
			55118: outdata = 32'd10418;
			55119: outdata = 32'd10417;
			55120: outdata = 32'd10416;
			55121: outdata = 32'd10415;
			55122: outdata = 32'd10414;
			55123: outdata = 32'd10413;
			55124: outdata = 32'd10412;
			55125: outdata = 32'd10411;
			55126: outdata = 32'd10410;
			55127: outdata = 32'd10409;
			55128: outdata = 32'd10408;
			55129: outdata = 32'd10407;
			55130: outdata = 32'd10406;
			55131: outdata = 32'd10405;
			55132: outdata = 32'd10404;
			55133: outdata = 32'd10403;
			55134: outdata = 32'd10402;
			55135: outdata = 32'd10401;
			55136: outdata = 32'd10400;
			55137: outdata = 32'd10399;
			55138: outdata = 32'd10398;
			55139: outdata = 32'd10397;
			55140: outdata = 32'd10396;
			55141: outdata = 32'd10395;
			55142: outdata = 32'd10394;
			55143: outdata = 32'd10393;
			55144: outdata = 32'd10392;
			55145: outdata = 32'd10391;
			55146: outdata = 32'd10390;
			55147: outdata = 32'd10389;
			55148: outdata = 32'd10388;
			55149: outdata = 32'd10387;
			55150: outdata = 32'd10386;
			55151: outdata = 32'd10385;
			55152: outdata = 32'd10384;
			55153: outdata = 32'd10383;
			55154: outdata = 32'd10382;
			55155: outdata = 32'd10381;
			55156: outdata = 32'd10380;
			55157: outdata = 32'd10379;
			55158: outdata = 32'd10378;
			55159: outdata = 32'd10377;
			55160: outdata = 32'd10376;
			55161: outdata = 32'd10375;
			55162: outdata = 32'd10374;
			55163: outdata = 32'd10373;
			55164: outdata = 32'd10372;
			55165: outdata = 32'd10371;
			55166: outdata = 32'd10370;
			55167: outdata = 32'd10369;
			55168: outdata = 32'd10368;
			55169: outdata = 32'd10367;
			55170: outdata = 32'd10366;
			55171: outdata = 32'd10365;
			55172: outdata = 32'd10364;
			55173: outdata = 32'd10363;
			55174: outdata = 32'd10362;
			55175: outdata = 32'd10361;
			55176: outdata = 32'd10360;
			55177: outdata = 32'd10359;
			55178: outdata = 32'd10358;
			55179: outdata = 32'd10357;
			55180: outdata = 32'd10356;
			55181: outdata = 32'd10355;
			55182: outdata = 32'd10354;
			55183: outdata = 32'd10353;
			55184: outdata = 32'd10352;
			55185: outdata = 32'd10351;
			55186: outdata = 32'd10350;
			55187: outdata = 32'd10349;
			55188: outdata = 32'd10348;
			55189: outdata = 32'd10347;
			55190: outdata = 32'd10346;
			55191: outdata = 32'd10345;
			55192: outdata = 32'd10344;
			55193: outdata = 32'd10343;
			55194: outdata = 32'd10342;
			55195: outdata = 32'd10341;
			55196: outdata = 32'd10340;
			55197: outdata = 32'd10339;
			55198: outdata = 32'd10338;
			55199: outdata = 32'd10337;
			55200: outdata = 32'd10336;
			55201: outdata = 32'd10335;
			55202: outdata = 32'd10334;
			55203: outdata = 32'd10333;
			55204: outdata = 32'd10332;
			55205: outdata = 32'd10331;
			55206: outdata = 32'd10330;
			55207: outdata = 32'd10329;
			55208: outdata = 32'd10328;
			55209: outdata = 32'd10327;
			55210: outdata = 32'd10326;
			55211: outdata = 32'd10325;
			55212: outdata = 32'd10324;
			55213: outdata = 32'd10323;
			55214: outdata = 32'd10322;
			55215: outdata = 32'd10321;
			55216: outdata = 32'd10320;
			55217: outdata = 32'd10319;
			55218: outdata = 32'd10318;
			55219: outdata = 32'd10317;
			55220: outdata = 32'd10316;
			55221: outdata = 32'd10315;
			55222: outdata = 32'd10314;
			55223: outdata = 32'd10313;
			55224: outdata = 32'd10312;
			55225: outdata = 32'd10311;
			55226: outdata = 32'd10310;
			55227: outdata = 32'd10309;
			55228: outdata = 32'd10308;
			55229: outdata = 32'd10307;
			55230: outdata = 32'd10306;
			55231: outdata = 32'd10305;
			55232: outdata = 32'd10304;
			55233: outdata = 32'd10303;
			55234: outdata = 32'd10302;
			55235: outdata = 32'd10301;
			55236: outdata = 32'd10300;
			55237: outdata = 32'd10299;
			55238: outdata = 32'd10298;
			55239: outdata = 32'd10297;
			55240: outdata = 32'd10296;
			55241: outdata = 32'd10295;
			55242: outdata = 32'd10294;
			55243: outdata = 32'd10293;
			55244: outdata = 32'd10292;
			55245: outdata = 32'd10291;
			55246: outdata = 32'd10290;
			55247: outdata = 32'd10289;
			55248: outdata = 32'd10288;
			55249: outdata = 32'd10287;
			55250: outdata = 32'd10286;
			55251: outdata = 32'd10285;
			55252: outdata = 32'd10284;
			55253: outdata = 32'd10283;
			55254: outdata = 32'd10282;
			55255: outdata = 32'd10281;
			55256: outdata = 32'd10280;
			55257: outdata = 32'd10279;
			55258: outdata = 32'd10278;
			55259: outdata = 32'd10277;
			55260: outdata = 32'd10276;
			55261: outdata = 32'd10275;
			55262: outdata = 32'd10274;
			55263: outdata = 32'd10273;
			55264: outdata = 32'd10272;
			55265: outdata = 32'd10271;
			55266: outdata = 32'd10270;
			55267: outdata = 32'd10269;
			55268: outdata = 32'd10268;
			55269: outdata = 32'd10267;
			55270: outdata = 32'd10266;
			55271: outdata = 32'd10265;
			55272: outdata = 32'd10264;
			55273: outdata = 32'd10263;
			55274: outdata = 32'd10262;
			55275: outdata = 32'd10261;
			55276: outdata = 32'd10260;
			55277: outdata = 32'd10259;
			55278: outdata = 32'd10258;
			55279: outdata = 32'd10257;
			55280: outdata = 32'd10256;
			55281: outdata = 32'd10255;
			55282: outdata = 32'd10254;
			55283: outdata = 32'd10253;
			55284: outdata = 32'd10252;
			55285: outdata = 32'd10251;
			55286: outdata = 32'd10250;
			55287: outdata = 32'd10249;
			55288: outdata = 32'd10248;
			55289: outdata = 32'd10247;
			55290: outdata = 32'd10246;
			55291: outdata = 32'd10245;
			55292: outdata = 32'd10244;
			55293: outdata = 32'd10243;
			55294: outdata = 32'd10242;
			55295: outdata = 32'd10241;
			55296: outdata = 32'd10240;
			55297: outdata = 32'd10239;
			55298: outdata = 32'd10238;
			55299: outdata = 32'd10237;
			55300: outdata = 32'd10236;
			55301: outdata = 32'd10235;
			55302: outdata = 32'd10234;
			55303: outdata = 32'd10233;
			55304: outdata = 32'd10232;
			55305: outdata = 32'd10231;
			55306: outdata = 32'd10230;
			55307: outdata = 32'd10229;
			55308: outdata = 32'd10228;
			55309: outdata = 32'd10227;
			55310: outdata = 32'd10226;
			55311: outdata = 32'd10225;
			55312: outdata = 32'd10224;
			55313: outdata = 32'd10223;
			55314: outdata = 32'd10222;
			55315: outdata = 32'd10221;
			55316: outdata = 32'd10220;
			55317: outdata = 32'd10219;
			55318: outdata = 32'd10218;
			55319: outdata = 32'd10217;
			55320: outdata = 32'd10216;
			55321: outdata = 32'd10215;
			55322: outdata = 32'd10214;
			55323: outdata = 32'd10213;
			55324: outdata = 32'd10212;
			55325: outdata = 32'd10211;
			55326: outdata = 32'd10210;
			55327: outdata = 32'd10209;
			55328: outdata = 32'd10208;
			55329: outdata = 32'd10207;
			55330: outdata = 32'd10206;
			55331: outdata = 32'd10205;
			55332: outdata = 32'd10204;
			55333: outdata = 32'd10203;
			55334: outdata = 32'd10202;
			55335: outdata = 32'd10201;
			55336: outdata = 32'd10200;
			55337: outdata = 32'd10199;
			55338: outdata = 32'd10198;
			55339: outdata = 32'd10197;
			55340: outdata = 32'd10196;
			55341: outdata = 32'd10195;
			55342: outdata = 32'd10194;
			55343: outdata = 32'd10193;
			55344: outdata = 32'd10192;
			55345: outdata = 32'd10191;
			55346: outdata = 32'd10190;
			55347: outdata = 32'd10189;
			55348: outdata = 32'd10188;
			55349: outdata = 32'd10187;
			55350: outdata = 32'd10186;
			55351: outdata = 32'd10185;
			55352: outdata = 32'd10184;
			55353: outdata = 32'd10183;
			55354: outdata = 32'd10182;
			55355: outdata = 32'd10181;
			55356: outdata = 32'd10180;
			55357: outdata = 32'd10179;
			55358: outdata = 32'd10178;
			55359: outdata = 32'd10177;
			55360: outdata = 32'd10176;
			55361: outdata = 32'd10175;
			55362: outdata = 32'd10174;
			55363: outdata = 32'd10173;
			55364: outdata = 32'd10172;
			55365: outdata = 32'd10171;
			55366: outdata = 32'd10170;
			55367: outdata = 32'd10169;
			55368: outdata = 32'd10168;
			55369: outdata = 32'd10167;
			55370: outdata = 32'd10166;
			55371: outdata = 32'd10165;
			55372: outdata = 32'd10164;
			55373: outdata = 32'd10163;
			55374: outdata = 32'd10162;
			55375: outdata = 32'd10161;
			55376: outdata = 32'd10160;
			55377: outdata = 32'd10159;
			55378: outdata = 32'd10158;
			55379: outdata = 32'd10157;
			55380: outdata = 32'd10156;
			55381: outdata = 32'd10155;
			55382: outdata = 32'd10154;
			55383: outdata = 32'd10153;
			55384: outdata = 32'd10152;
			55385: outdata = 32'd10151;
			55386: outdata = 32'd10150;
			55387: outdata = 32'd10149;
			55388: outdata = 32'd10148;
			55389: outdata = 32'd10147;
			55390: outdata = 32'd10146;
			55391: outdata = 32'd10145;
			55392: outdata = 32'd10144;
			55393: outdata = 32'd10143;
			55394: outdata = 32'd10142;
			55395: outdata = 32'd10141;
			55396: outdata = 32'd10140;
			55397: outdata = 32'd10139;
			55398: outdata = 32'd10138;
			55399: outdata = 32'd10137;
			55400: outdata = 32'd10136;
			55401: outdata = 32'd10135;
			55402: outdata = 32'd10134;
			55403: outdata = 32'd10133;
			55404: outdata = 32'd10132;
			55405: outdata = 32'd10131;
			55406: outdata = 32'd10130;
			55407: outdata = 32'd10129;
			55408: outdata = 32'd10128;
			55409: outdata = 32'd10127;
			55410: outdata = 32'd10126;
			55411: outdata = 32'd10125;
			55412: outdata = 32'd10124;
			55413: outdata = 32'd10123;
			55414: outdata = 32'd10122;
			55415: outdata = 32'd10121;
			55416: outdata = 32'd10120;
			55417: outdata = 32'd10119;
			55418: outdata = 32'd10118;
			55419: outdata = 32'd10117;
			55420: outdata = 32'd10116;
			55421: outdata = 32'd10115;
			55422: outdata = 32'd10114;
			55423: outdata = 32'd10113;
			55424: outdata = 32'd10112;
			55425: outdata = 32'd10111;
			55426: outdata = 32'd10110;
			55427: outdata = 32'd10109;
			55428: outdata = 32'd10108;
			55429: outdata = 32'd10107;
			55430: outdata = 32'd10106;
			55431: outdata = 32'd10105;
			55432: outdata = 32'd10104;
			55433: outdata = 32'd10103;
			55434: outdata = 32'd10102;
			55435: outdata = 32'd10101;
			55436: outdata = 32'd10100;
			55437: outdata = 32'd10099;
			55438: outdata = 32'd10098;
			55439: outdata = 32'd10097;
			55440: outdata = 32'd10096;
			55441: outdata = 32'd10095;
			55442: outdata = 32'd10094;
			55443: outdata = 32'd10093;
			55444: outdata = 32'd10092;
			55445: outdata = 32'd10091;
			55446: outdata = 32'd10090;
			55447: outdata = 32'd10089;
			55448: outdata = 32'd10088;
			55449: outdata = 32'd10087;
			55450: outdata = 32'd10086;
			55451: outdata = 32'd10085;
			55452: outdata = 32'd10084;
			55453: outdata = 32'd10083;
			55454: outdata = 32'd10082;
			55455: outdata = 32'd10081;
			55456: outdata = 32'd10080;
			55457: outdata = 32'd10079;
			55458: outdata = 32'd10078;
			55459: outdata = 32'd10077;
			55460: outdata = 32'd10076;
			55461: outdata = 32'd10075;
			55462: outdata = 32'd10074;
			55463: outdata = 32'd10073;
			55464: outdata = 32'd10072;
			55465: outdata = 32'd10071;
			55466: outdata = 32'd10070;
			55467: outdata = 32'd10069;
			55468: outdata = 32'd10068;
			55469: outdata = 32'd10067;
			55470: outdata = 32'd10066;
			55471: outdata = 32'd10065;
			55472: outdata = 32'd10064;
			55473: outdata = 32'd10063;
			55474: outdata = 32'd10062;
			55475: outdata = 32'd10061;
			55476: outdata = 32'd10060;
			55477: outdata = 32'd10059;
			55478: outdata = 32'd10058;
			55479: outdata = 32'd10057;
			55480: outdata = 32'd10056;
			55481: outdata = 32'd10055;
			55482: outdata = 32'd10054;
			55483: outdata = 32'd10053;
			55484: outdata = 32'd10052;
			55485: outdata = 32'd10051;
			55486: outdata = 32'd10050;
			55487: outdata = 32'd10049;
			55488: outdata = 32'd10048;
			55489: outdata = 32'd10047;
			55490: outdata = 32'd10046;
			55491: outdata = 32'd10045;
			55492: outdata = 32'd10044;
			55493: outdata = 32'd10043;
			55494: outdata = 32'd10042;
			55495: outdata = 32'd10041;
			55496: outdata = 32'd10040;
			55497: outdata = 32'd10039;
			55498: outdata = 32'd10038;
			55499: outdata = 32'd10037;
			55500: outdata = 32'd10036;
			55501: outdata = 32'd10035;
			55502: outdata = 32'd10034;
			55503: outdata = 32'd10033;
			55504: outdata = 32'd10032;
			55505: outdata = 32'd10031;
			55506: outdata = 32'd10030;
			55507: outdata = 32'd10029;
			55508: outdata = 32'd10028;
			55509: outdata = 32'd10027;
			55510: outdata = 32'd10026;
			55511: outdata = 32'd10025;
			55512: outdata = 32'd10024;
			55513: outdata = 32'd10023;
			55514: outdata = 32'd10022;
			55515: outdata = 32'd10021;
			55516: outdata = 32'd10020;
			55517: outdata = 32'd10019;
			55518: outdata = 32'd10018;
			55519: outdata = 32'd10017;
			55520: outdata = 32'd10016;
			55521: outdata = 32'd10015;
			55522: outdata = 32'd10014;
			55523: outdata = 32'd10013;
			55524: outdata = 32'd10012;
			55525: outdata = 32'd10011;
			55526: outdata = 32'd10010;
			55527: outdata = 32'd10009;
			55528: outdata = 32'd10008;
			55529: outdata = 32'd10007;
			55530: outdata = 32'd10006;
			55531: outdata = 32'd10005;
			55532: outdata = 32'd10004;
			55533: outdata = 32'd10003;
			55534: outdata = 32'd10002;
			55535: outdata = 32'd10001;
			55536: outdata = 32'd10000;
			55537: outdata = 32'd9999;
			55538: outdata = 32'd9998;
			55539: outdata = 32'd9997;
			55540: outdata = 32'd9996;
			55541: outdata = 32'd9995;
			55542: outdata = 32'd9994;
			55543: outdata = 32'd9993;
			55544: outdata = 32'd9992;
			55545: outdata = 32'd9991;
			55546: outdata = 32'd9990;
			55547: outdata = 32'd9989;
			55548: outdata = 32'd9988;
			55549: outdata = 32'd9987;
			55550: outdata = 32'd9986;
			55551: outdata = 32'd9985;
			55552: outdata = 32'd9984;
			55553: outdata = 32'd9983;
			55554: outdata = 32'd9982;
			55555: outdata = 32'd9981;
			55556: outdata = 32'd9980;
			55557: outdata = 32'd9979;
			55558: outdata = 32'd9978;
			55559: outdata = 32'd9977;
			55560: outdata = 32'd9976;
			55561: outdata = 32'd9975;
			55562: outdata = 32'd9974;
			55563: outdata = 32'd9973;
			55564: outdata = 32'd9972;
			55565: outdata = 32'd9971;
			55566: outdata = 32'd9970;
			55567: outdata = 32'd9969;
			55568: outdata = 32'd9968;
			55569: outdata = 32'd9967;
			55570: outdata = 32'd9966;
			55571: outdata = 32'd9965;
			55572: outdata = 32'd9964;
			55573: outdata = 32'd9963;
			55574: outdata = 32'd9962;
			55575: outdata = 32'd9961;
			55576: outdata = 32'd9960;
			55577: outdata = 32'd9959;
			55578: outdata = 32'd9958;
			55579: outdata = 32'd9957;
			55580: outdata = 32'd9956;
			55581: outdata = 32'd9955;
			55582: outdata = 32'd9954;
			55583: outdata = 32'd9953;
			55584: outdata = 32'd9952;
			55585: outdata = 32'd9951;
			55586: outdata = 32'd9950;
			55587: outdata = 32'd9949;
			55588: outdata = 32'd9948;
			55589: outdata = 32'd9947;
			55590: outdata = 32'd9946;
			55591: outdata = 32'd9945;
			55592: outdata = 32'd9944;
			55593: outdata = 32'd9943;
			55594: outdata = 32'd9942;
			55595: outdata = 32'd9941;
			55596: outdata = 32'd9940;
			55597: outdata = 32'd9939;
			55598: outdata = 32'd9938;
			55599: outdata = 32'd9937;
			55600: outdata = 32'd9936;
			55601: outdata = 32'd9935;
			55602: outdata = 32'd9934;
			55603: outdata = 32'd9933;
			55604: outdata = 32'd9932;
			55605: outdata = 32'd9931;
			55606: outdata = 32'd9930;
			55607: outdata = 32'd9929;
			55608: outdata = 32'd9928;
			55609: outdata = 32'd9927;
			55610: outdata = 32'd9926;
			55611: outdata = 32'd9925;
			55612: outdata = 32'd9924;
			55613: outdata = 32'd9923;
			55614: outdata = 32'd9922;
			55615: outdata = 32'd9921;
			55616: outdata = 32'd9920;
			55617: outdata = 32'd9919;
			55618: outdata = 32'd9918;
			55619: outdata = 32'd9917;
			55620: outdata = 32'd9916;
			55621: outdata = 32'd9915;
			55622: outdata = 32'd9914;
			55623: outdata = 32'd9913;
			55624: outdata = 32'd9912;
			55625: outdata = 32'd9911;
			55626: outdata = 32'd9910;
			55627: outdata = 32'd9909;
			55628: outdata = 32'd9908;
			55629: outdata = 32'd9907;
			55630: outdata = 32'd9906;
			55631: outdata = 32'd9905;
			55632: outdata = 32'd9904;
			55633: outdata = 32'd9903;
			55634: outdata = 32'd9902;
			55635: outdata = 32'd9901;
			55636: outdata = 32'd9900;
			55637: outdata = 32'd9899;
			55638: outdata = 32'd9898;
			55639: outdata = 32'd9897;
			55640: outdata = 32'd9896;
			55641: outdata = 32'd9895;
			55642: outdata = 32'd9894;
			55643: outdata = 32'd9893;
			55644: outdata = 32'd9892;
			55645: outdata = 32'd9891;
			55646: outdata = 32'd9890;
			55647: outdata = 32'd9889;
			55648: outdata = 32'd9888;
			55649: outdata = 32'd9887;
			55650: outdata = 32'd9886;
			55651: outdata = 32'd9885;
			55652: outdata = 32'd9884;
			55653: outdata = 32'd9883;
			55654: outdata = 32'd9882;
			55655: outdata = 32'd9881;
			55656: outdata = 32'd9880;
			55657: outdata = 32'd9879;
			55658: outdata = 32'd9878;
			55659: outdata = 32'd9877;
			55660: outdata = 32'd9876;
			55661: outdata = 32'd9875;
			55662: outdata = 32'd9874;
			55663: outdata = 32'd9873;
			55664: outdata = 32'd9872;
			55665: outdata = 32'd9871;
			55666: outdata = 32'd9870;
			55667: outdata = 32'd9869;
			55668: outdata = 32'd9868;
			55669: outdata = 32'd9867;
			55670: outdata = 32'd9866;
			55671: outdata = 32'd9865;
			55672: outdata = 32'd9864;
			55673: outdata = 32'd9863;
			55674: outdata = 32'd9862;
			55675: outdata = 32'd9861;
			55676: outdata = 32'd9860;
			55677: outdata = 32'd9859;
			55678: outdata = 32'd9858;
			55679: outdata = 32'd9857;
			55680: outdata = 32'd9856;
			55681: outdata = 32'd9855;
			55682: outdata = 32'd9854;
			55683: outdata = 32'd9853;
			55684: outdata = 32'd9852;
			55685: outdata = 32'd9851;
			55686: outdata = 32'd9850;
			55687: outdata = 32'd9849;
			55688: outdata = 32'd9848;
			55689: outdata = 32'd9847;
			55690: outdata = 32'd9846;
			55691: outdata = 32'd9845;
			55692: outdata = 32'd9844;
			55693: outdata = 32'd9843;
			55694: outdata = 32'd9842;
			55695: outdata = 32'd9841;
			55696: outdata = 32'd9840;
			55697: outdata = 32'd9839;
			55698: outdata = 32'd9838;
			55699: outdata = 32'd9837;
			55700: outdata = 32'd9836;
			55701: outdata = 32'd9835;
			55702: outdata = 32'd9834;
			55703: outdata = 32'd9833;
			55704: outdata = 32'd9832;
			55705: outdata = 32'd9831;
			55706: outdata = 32'd9830;
			55707: outdata = 32'd9829;
			55708: outdata = 32'd9828;
			55709: outdata = 32'd9827;
			55710: outdata = 32'd9826;
			55711: outdata = 32'd9825;
			55712: outdata = 32'd9824;
			55713: outdata = 32'd9823;
			55714: outdata = 32'd9822;
			55715: outdata = 32'd9821;
			55716: outdata = 32'd9820;
			55717: outdata = 32'd9819;
			55718: outdata = 32'd9818;
			55719: outdata = 32'd9817;
			55720: outdata = 32'd9816;
			55721: outdata = 32'd9815;
			55722: outdata = 32'd9814;
			55723: outdata = 32'd9813;
			55724: outdata = 32'd9812;
			55725: outdata = 32'd9811;
			55726: outdata = 32'd9810;
			55727: outdata = 32'd9809;
			55728: outdata = 32'd9808;
			55729: outdata = 32'd9807;
			55730: outdata = 32'd9806;
			55731: outdata = 32'd9805;
			55732: outdata = 32'd9804;
			55733: outdata = 32'd9803;
			55734: outdata = 32'd9802;
			55735: outdata = 32'd9801;
			55736: outdata = 32'd9800;
			55737: outdata = 32'd9799;
			55738: outdata = 32'd9798;
			55739: outdata = 32'd9797;
			55740: outdata = 32'd9796;
			55741: outdata = 32'd9795;
			55742: outdata = 32'd9794;
			55743: outdata = 32'd9793;
			55744: outdata = 32'd9792;
			55745: outdata = 32'd9791;
			55746: outdata = 32'd9790;
			55747: outdata = 32'd9789;
			55748: outdata = 32'd9788;
			55749: outdata = 32'd9787;
			55750: outdata = 32'd9786;
			55751: outdata = 32'd9785;
			55752: outdata = 32'd9784;
			55753: outdata = 32'd9783;
			55754: outdata = 32'd9782;
			55755: outdata = 32'd9781;
			55756: outdata = 32'd9780;
			55757: outdata = 32'd9779;
			55758: outdata = 32'd9778;
			55759: outdata = 32'd9777;
			55760: outdata = 32'd9776;
			55761: outdata = 32'd9775;
			55762: outdata = 32'd9774;
			55763: outdata = 32'd9773;
			55764: outdata = 32'd9772;
			55765: outdata = 32'd9771;
			55766: outdata = 32'd9770;
			55767: outdata = 32'd9769;
			55768: outdata = 32'd9768;
			55769: outdata = 32'd9767;
			55770: outdata = 32'd9766;
			55771: outdata = 32'd9765;
			55772: outdata = 32'd9764;
			55773: outdata = 32'd9763;
			55774: outdata = 32'd9762;
			55775: outdata = 32'd9761;
			55776: outdata = 32'd9760;
			55777: outdata = 32'd9759;
			55778: outdata = 32'd9758;
			55779: outdata = 32'd9757;
			55780: outdata = 32'd9756;
			55781: outdata = 32'd9755;
			55782: outdata = 32'd9754;
			55783: outdata = 32'd9753;
			55784: outdata = 32'd9752;
			55785: outdata = 32'd9751;
			55786: outdata = 32'd9750;
			55787: outdata = 32'd9749;
			55788: outdata = 32'd9748;
			55789: outdata = 32'd9747;
			55790: outdata = 32'd9746;
			55791: outdata = 32'd9745;
			55792: outdata = 32'd9744;
			55793: outdata = 32'd9743;
			55794: outdata = 32'd9742;
			55795: outdata = 32'd9741;
			55796: outdata = 32'd9740;
			55797: outdata = 32'd9739;
			55798: outdata = 32'd9738;
			55799: outdata = 32'd9737;
			55800: outdata = 32'd9736;
			55801: outdata = 32'd9735;
			55802: outdata = 32'd9734;
			55803: outdata = 32'd9733;
			55804: outdata = 32'd9732;
			55805: outdata = 32'd9731;
			55806: outdata = 32'd9730;
			55807: outdata = 32'd9729;
			55808: outdata = 32'd9728;
			55809: outdata = 32'd9727;
			55810: outdata = 32'd9726;
			55811: outdata = 32'd9725;
			55812: outdata = 32'd9724;
			55813: outdata = 32'd9723;
			55814: outdata = 32'd9722;
			55815: outdata = 32'd9721;
			55816: outdata = 32'd9720;
			55817: outdata = 32'd9719;
			55818: outdata = 32'd9718;
			55819: outdata = 32'd9717;
			55820: outdata = 32'd9716;
			55821: outdata = 32'd9715;
			55822: outdata = 32'd9714;
			55823: outdata = 32'd9713;
			55824: outdata = 32'd9712;
			55825: outdata = 32'd9711;
			55826: outdata = 32'd9710;
			55827: outdata = 32'd9709;
			55828: outdata = 32'd9708;
			55829: outdata = 32'd9707;
			55830: outdata = 32'd9706;
			55831: outdata = 32'd9705;
			55832: outdata = 32'd9704;
			55833: outdata = 32'd9703;
			55834: outdata = 32'd9702;
			55835: outdata = 32'd9701;
			55836: outdata = 32'd9700;
			55837: outdata = 32'd9699;
			55838: outdata = 32'd9698;
			55839: outdata = 32'd9697;
			55840: outdata = 32'd9696;
			55841: outdata = 32'd9695;
			55842: outdata = 32'd9694;
			55843: outdata = 32'd9693;
			55844: outdata = 32'd9692;
			55845: outdata = 32'd9691;
			55846: outdata = 32'd9690;
			55847: outdata = 32'd9689;
			55848: outdata = 32'd9688;
			55849: outdata = 32'd9687;
			55850: outdata = 32'd9686;
			55851: outdata = 32'd9685;
			55852: outdata = 32'd9684;
			55853: outdata = 32'd9683;
			55854: outdata = 32'd9682;
			55855: outdata = 32'd9681;
			55856: outdata = 32'd9680;
			55857: outdata = 32'd9679;
			55858: outdata = 32'd9678;
			55859: outdata = 32'd9677;
			55860: outdata = 32'd9676;
			55861: outdata = 32'd9675;
			55862: outdata = 32'd9674;
			55863: outdata = 32'd9673;
			55864: outdata = 32'd9672;
			55865: outdata = 32'd9671;
			55866: outdata = 32'd9670;
			55867: outdata = 32'd9669;
			55868: outdata = 32'd9668;
			55869: outdata = 32'd9667;
			55870: outdata = 32'd9666;
			55871: outdata = 32'd9665;
			55872: outdata = 32'd9664;
			55873: outdata = 32'd9663;
			55874: outdata = 32'd9662;
			55875: outdata = 32'd9661;
			55876: outdata = 32'd9660;
			55877: outdata = 32'd9659;
			55878: outdata = 32'd9658;
			55879: outdata = 32'd9657;
			55880: outdata = 32'd9656;
			55881: outdata = 32'd9655;
			55882: outdata = 32'd9654;
			55883: outdata = 32'd9653;
			55884: outdata = 32'd9652;
			55885: outdata = 32'd9651;
			55886: outdata = 32'd9650;
			55887: outdata = 32'd9649;
			55888: outdata = 32'd9648;
			55889: outdata = 32'd9647;
			55890: outdata = 32'd9646;
			55891: outdata = 32'd9645;
			55892: outdata = 32'd9644;
			55893: outdata = 32'd9643;
			55894: outdata = 32'd9642;
			55895: outdata = 32'd9641;
			55896: outdata = 32'd9640;
			55897: outdata = 32'd9639;
			55898: outdata = 32'd9638;
			55899: outdata = 32'd9637;
			55900: outdata = 32'd9636;
			55901: outdata = 32'd9635;
			55902: outdata = 32'd9634;
			55903: outdata = 32'd9633;
			55904: outdata = 32'd9632;
			55905: outdata = 32'd9631;
			55906: outdata = 32'd9630;
			55907: outdata = 32'd9629;
			55908: outdata = 32'd9628;
			55909: outdata = 32'd9627;
			55910: outdata = 32'd9626;
			55911: outdata = 32'd9625;
			55912: outdata = 32'd9624;
			55913: outdata = 32'd9623;
			55914: outdata = 32'd9622;
			55915: outdata = 32'd9621;
			55916: outdata = 32'd9620;
			55917: outdata = 32'd9619;
			55918: outdata = 32'd9618;
			55919: outdata = 32'd9617;
			55920: outdata = 32'd9616;
			55921: outdata = 32'd9615;
			55922: outdata = 32'd9614;
			55923: outdata = 32'd9613;
			55924: outdata = 32'd9612;
			55925: outdata = 32'd9611;
			55926: outdata = 32'd9610;
			55927: outdata = 32'd9609;
			55928: outdata = 32'd9608;
			55929: outdata = 32'd9607;
			55930: outdata = 32'd9606;
			55931: outdata = 32'd9605;
			55932: outdata = 32'd9604;
			55933: outdata = 32'd9603;
			55934: outdata = 32'd9602;
			55935: outdata = 32'd9601;
			55936: outdata = 32'd9600;
			55937: outdata = 32'd9599;
			55938: outdata = 32'd9598;
			55939: outdata = 32'd9597;
			55940: outdata = 32'd9596;
			55941: outdata = 32'd9595;
			55942: outdata = 32'd9594;
			55943: outdata = 32'd9593;
			55944: outdata = 32'd9592;
			55945: outdata = 32'd9591;
			55946: outdata = 32'd9590;
			55947: outdata = 32'd9589;
			55948: outdata = 32'd9588;
			55949: outdata = 32'd9587;
			55950: outdata = 32'd9586;
			55951: outdata = 32'd9585;
			55952: outdata = 32'd9584;
			55953: outdata = 32'd9583;
			55954: outdata = 32'd9582;
			55955: outdata = 32'd9581;
			55956: outdata = 32'd9580;
			55957: outdata = 32'd9579;
			55958: outdata = 32'd9578;
			55959: outdata = 32'd9577;
			55960: outdata = 32'd9576;
			55961: outdata = 32'd9575;
			55962: outdata = 32'd9574;
			55963: outdata = 32'd9573;
			55964: outdata = 32'd9572;
			55965: outdata = 32'd9571;
			55966: outdata = 32'd9570;
			55967: outdata = 32'd9569;
			55968: outdata = 32'd9568;
			55969: outdata = 32'd9567;
			55970: outdata = 32'd9566;
			55971: outdata = 32'd9565;
			55972: outdata = 32'd9564;
			55973: outdata = 32'd9563;
			55974: outdata = 32'd9562;
			55975: outdata = 32'd9561;
			55976: outdata = 32'd9560;
			55977: outdata = 32'd9559;
			55978: outdata = 32'd9558;
			55979: outdata = 32'd9557;
			55980: outdata = 32'd9556;
			55981: outdata = 32'd9555;
			55982: outdata = 32'd9554;
			55983: outdata = 32'd9553;
			55984: outdata = 32'd9552;
			55985: outdata = 32'd9551;
			55986: outdata = 32'd9550;
			55987: outdata = 32'd9549;
			55988: outdata = 32'd9548;
			55989: outdata = 32'd9547;
			55990: outdata = 32'd9546;
			55991: outdata = 32'd9545;
			55992: outdata = 32'd9544;
			55993: outdata = 32'd9543;
			55994: outdata = 32'd9542;
			55995: outdata = 32'd9541;
			55996: outdata = 32'd9540;
			55997: outdata = 32'd9539;
			55998: outdata = 32'd9538;
			55999: outdata = 32'd9537;
			56000: outdata = 32'd9536;
			56001: outdata = 32'd9535;
			56002: outdata = 32'd9534;
			56003: outdata = 32'd9533;
			56004: outdata = 32'd9532;
			56005: outdata = 32'd9531;
			56006: outdata = 32'd9530;
			56007: outdata = 32'd9529;
			56008: outdata = 32'd9528;
			56009: outdata = 32'd9527;
			56010: outdata = 32'd9526;
			56011: outdata = 32'd9525;
			56012: outdata = 32'd9524;
			56013: outdata = 32'd9523;
			56014: outdata = 32'd9522;
			56015: outdata = 32'd9521;
			56016: outdata = 32'd9520;
			56017: outdata = 32'd9519;
			56018: outdata = 32'd9518;
			56019: outdata = 32'd9517;
			56020: outdata = 32'd9516;
			56021: outdata = 32'd9515;
			56022: outdata = 32'd9514;
			56023: outdata = 32'd9513;
			56024: outdata = 32'd9512;
			56025: outdata = 32'd9511;
			56026: outdata = 32'd9510;
			56027: outdata = 32'd9509;
			56028: outdata = 32'd9508;
			56029: outdata = 32'd9507;
			56030: outdata = 32'd9506;
			56031: outdata = 32'd9505;
			56032: outdata = 32'd9504;
			56033: outdata = 32'd9503;
			56034: outdata = 32'd9502;
			56035: outdata = 32'd9501;
			56036: outdata = 32'd9500;
			56037: outdata = 32'd9499;
			56038: outdata = 32'd9498;
			56039: outdata = 32'd9497;
			56040: outdata = 32'd9496;
			56041: outdata = 32'd9495;
			56042: outdata = 32'd9494;
			56043: outdata = 32'd9493;
			56044: outdata = 32'd9492;
			56045: outdata = 32'd9491;
			56046: outdata = 32'd9490;
			56047: outdata = 32'd9489;
			56048: outdata = 32'd9488;
			56049: outdata = 32'd9487;
			56050: outdata = 32'd9486;
			56051: outdata = 32'd9485;
			56052: outdata = 32'd9484;
			56053: outdata = 32'd9483;
			56054: outdata = 32'd9482;
			56055: outdata = 32'd9481;
			56056: outdata = 32'd9480;
			56057: outdata = 32'd9479;
			56058: outdata = 32'd9478;
			56059: outdata = 32'd9477;
			56060: outdata = 32'd9476;
			56061: outdata = 32'd9475;
			56062: outdata = 32'd9474;
			56063: outdata = 32'd9473;
			56064: outdata = 32'd9472;
			56065: outdata = 32'd9471;
			56066: outdata = 32'd9470;
			56067: outdata = 32'd9469;
			56068: outdata = 32'd9468;
			56069: outdata = 32'd9467;
			56070: outdata = 32'd9466;
			56071: outdata = 32'd9465;
			56072: outdata = 32'd9464;
			56073: outdata = 32'd9463;
			56074: outdata = 32'd9462;
			56075: outdata = 32'd9461;
			56076: outdata = 32'd9460;
			56077: outdata = 32'd9459;
			56078: outdata = 32'd9458;
			56079: outdata = 32'd9457;
			56080: outdata = 32'd9456;
			56081: outdata = 32'd9455;
			56082: outdata = 32'd9454;
			56083: outdata = 32'd9453;
			56084: outdata = 32'd9452;
			56085: outdata = 32'd9451;
			56086: outdata = 32'd9450;
			56087: outdata = 32'd9449;
			56088: outdata = 32'd9448;
			56089: outdata = 32'd9447;
			56090: outdata = 32'd9446;
			56091: outdata = 32'd9445;
			56092: outdata = 32'd9444;
			56093: outdata = 32'd9443;
			56094: outdata = 32'd9442;
			56095: outdata = 32'd9441;
			56096: outdata = 32'd9440;
			56097: outdata = 32'd9439;
			56098: outdata = 32'd9438;
			56099: outdata = 32'd9437;
			56100: outdata = 32'd9436;
			56101: outdata = 32'd9435;
			56102: outdata = 32'd9434;
			56103: outdata = 32'd9433;
			56104: outdata = 32'd9432;
			56105: outdata = 32'd9431;
			56106: outdata = 32'd9430;
			56107: outdata = 32'd9429;
			56108: outdata = 32'd9428;
			56109: outdata = 32'd9427;
			56110: outdata = 32'd9426;
			56111: outdata = 32'd9425;
			56112: outdata = 32'd9424;
			56113: outdata = 32'd9423;
			56114: outdata = 32'd9422;
			56115: outdata = 32'd9421;
			56116: outdata = 32'd9420;
			56117: outdata = 32'd9419;
			56118: outdata = 32'd9418;
			56119: outdata = 32'd9417;
			56120: outdata = 32'd9416;
			56121: outdata = 32'd9415;
			56122: outdata = 32'd9414;
			56123: outdata = 32'd9413;
			56124: outdata = 32'd9412;
			56125: outdata = 32'd9411;
			56126: outdata = 32'd9410;
			56127: outdata = 32'd9409;
			56128: outdata = 32'd9408;
			56129: outdata = 32'd9407;
			56130: outdata = 32'd9406;
			56131: outdata = 32'd9405;
			56132: outdata = 32'd9404;
			56133: outdata = 32'd9403;
			56134: outdata = 32'd9402;
			56135: outdata = 32'd9401;
			56136: outdata = 32'd9400;
			56137: outdata = 32'd9399;
			56138: outdata = 32'd9398;
			56139: outdata = 32'd9397;
			56140: outdata = 32'd9396;
			56141: outdata = 32'd9395;
			56142: outdata = 32'd9394;
			56143: outdata = 32'd9393;
			56144: outdata = 32'd9392;
			56145: outdata = 32'd9391;
			56146: outdata = 32'd9390;
			56147: outdata = 32'd9389;
			56148: outdata = 32'd9388;
			56149: outdata = 32'd9387;
			56150: outdata = 32'd9386;
			56151: outdata = 32'd9385;
			56152: outdata = 32'd9384;
			56153: outdata = 32'd9383;
			56154: outdata = 32'd9382;
			56155: outdata = 32'd9381;
			56156: outdata = 32'd9380;
			56157: outdata = 32'd9379;
			56158: outdata = 32'd9378;
			56159: outdata = 32'd9377;
			56160: outdata = 32'd9376;
			56161: outdata = 32'd9375;
			56162: outdata = 32'd9374;
			56163: outdata = 32'd9373;
			56164: outdata = 32'd9372;
			56165: outdata = 32'd9371;
			56166: outdata = 32'd9370;
			56167: outdata = 32'd9369;
			56168: outdata = 32'd9368;
			56169: outdata = 32'd9367;
			56170: outdata = 32'd9366;
			56171: outdata = 32'd9365;
			56172: outdata = 32'd9364;
			56173: outdata = 32'd9363;
			56174: outdata = 32'd9362;
			56175: outdata = 32'd9361;
			56176: outdata = 32'd9360;
			56177: outdata = 32'd9359;
			56178: outdata = 32'd9358;
			56179: outdata = 32'd9357;
			56180: outdata = 32'd9356;
			56181: outdata = 32'd9355;
			56182: outdata = 32'd9354;
			56183: outdata = 32'd9353;
			56184: outdata = 32'd9352;
			56185: outdata = 32'd9351;
			56186: outdata = 32'd9350;
			56187: outdata = 32'd9349;
			56188: outdata = 32'd9348;
			56189: outdata = 32'd9347;
			56190: outdata = 32'd9346;
			56191: outdata = 32'd9345;
			56192: outdata = 32'd9344;
			56193: outdata = 32'd9343;
			56194: outdata = 32'd9342;
			56195: outdata = 32'd9341;
			56196: outdata = 32'd9340;
			56197: outdata = 32'd9339;
			56198: outdata = 32'd9338;
			56199: outdata = 32'd9337;
			56200: outdata = 32'd9336;
			56201: outdata = 32'd9335;
			56202: outdata = 32'd9334;
			56203: outdata = 32'd9333;
			56204: outdata = 32'd9332;
			56205: outdata = 32'd9331;
			56206: outdata = 32'd9330;
			56207: outdata = 32'd9329;
			56208: outdata = 32'd9328;
			56209: outdata = 32'd9327;
			56210: outdata = 32'd9326;
			56211: outdata = 32'd9325;
			56212: outdata = 32'd9324;
			56213: outdata = 32'd9323;
			56214: outdata = 32'd9322;
			56215: outdata = 32'd9321;
			56216: outdata = 32'd9320;
			56217: outdata = 32'd9319;
			56218: outdata = 32'd9318;
			56219: outdata = 32'd9317;
			56220: outdata = 32'd9316;
			56221: outdata = 32'd9315;
			56222: outdata = 32'd9314;
			56223: outdata = 32'd9313;
			56224: outdata = 32'd9312;
			56225: outdata = 32'd9311;
			56226: outdata = 32'd9310;
			56227: outdata = 32'd9309;
			56228: outdata = 32'd9308;
			56229: outdata = 32'd9307;
			56230: outdata = 32'd9306;
			56231: outdata = 32'd9305;
			56232: outdata = 32'd9304;
			56233: outdata = 32'd9303;
			56234: outdata = 32'd9302;
			56235: outdata = 32'd9301;
			56236: outdata = 32'd9300;
			56237: outdata = 32'd9299;
			56238: outdata = 32'd9298;
			56239: outdata = 32'd9297;
			56240: outdata = 32'd9296;
			56241: outdata = 32'd9295;
			56242: outdata = 32'd9294;
			56243: outdata = 32'd9293;
			56244: outdata = 32'd9292;
			56245: outdata = 32'd9291;
			56246: outdata = 32'd9290;
			56247: outdata = 32'd9289;
			56248: outdata = 32'd9288;
			56249: outdata = 32'd9287;
			56250: outdata = 32'd9286;
			56251: outdata = 32'd9285;
			56252: outdata = 32'd9284;
			56253: outdata = 32'd9283;
			56254: outdata = 32'd9282;
			56255: outdata = 32'd9281;
			56256: outdata = 32'd9280;
			56257: outdata = 32'd9279;
			56258: outdata = 32'd9278;
			56259: outdata = 32'd9277;
			56260: outdata = 32'd9276;
			56261: outdata = 32'd9275;
			56262: outdata = 32'd9274;
			56263: outdata = 32'd9273;
			56264: outdata = 32'd9272;
			56265: outdata = 32'd9271;
			56266: outdata = 32'd9270;
			56267: outdata = 32'd9269;
			56268: outdata = 32'd9268;
			56269: outdata = 32'd9267;
			56270: outdata = 32'd9266;
			56271: outdata = 32'd9265;
			56272: outdata = 32'd9264;
			56273: outdata = 32'd9263;
			56274: outdata = 32'd9262;
			56275: outdata = 32'd9261;
			56276: outdata = 32'd9260;
			56277: outdata = 32'd9259;
			56278: outdata = 32'd9258;
			56279: outdata = 32'd9257;
			56280: outdata = 32'd9256;
			56281: outdata = 32'd9255;
			56282: outdata = 32'd9254;
			56283: outdata = 32'd9253;
			56284: outdata = 32'd9252;
			56285: outdata = 32'd9251;
			56286: outdata = 32'd9250;
			56287: outdata = 32'd9249;
			56288: outdata = 32'd9248;
			56289: outdata = 32'd9247;
			56290: outdata = 32'd9246;
			56291: outdata = 32'd9245;
			56292: outdata = 32'd9244;
			56293: outdata = 32'd9243;
			56294: outdata = 32'd9242;
			56295: outdata = 32'd9241;
			56296: outdata = 32'd9240;
			56297: outdata = 32'd9239;
			56298: outdata = 32'd9238;
			56299: outdata = 32'd9237;
			56300: outdata = 32'd9236;
			56301: outdata = 32'd9235;
			56302: outdata = 32'd9234;
			56303: outdata = 32'd9233;
			56304: outdata = 32'd9232;
			56305: outdata = 32'd9231;
			56306: outdata = 32'd9230;
			56307: outdata = 32'd9229;
			56308: outdata = 32'd9228;
			56309: outdata = 32'd9227;
			56310: outdata = 32'd9226;
			56311: outdata = 32'd9225;
			56312: outdata = 32'd9224;
			56313: outdata = 32'd9223;
			56314: outdata = 32'd9222;
			56315: outdata = 32'd9221;
			56316: outdata = 32'd9220;
			56317: outdata = 32'd9219;
			56318: outdata = 32'd9218;
			56319: outdata = 32'd9217;
			56320: outdata = 32'd9216;
			56321: outdata = 32'd9215;
			56322: outdata = 32'd9214;
			56323: outdata = 32'd9213;
			56324: outdata = 32'd9212;
			56325: outdata = 32'd9211;
			56326: outdata = 32'd9210;
			56327: outdata = 32'd9209;
			56328: outdata = 32'd9208;
			56329: outdata = 32'd9207;
			56330: outdata = 32'd9206;
			56331: outdata = 32'd9205;
			56332: outdata = 32'd9204;
			56333: outdata = 32'd9203;
			56334: outdata = 32'd9202;
			56335: outdata = 32'd9201;
			56336: outdata = 32'd9200;
			56337: outdata = 32'd9199;
			56338: outdata = 32'd9198;
			56339: outdata = 32'd9197;
			56340: outdata = 32'd9196;
			56341: outdata = 32'd9195;
			56342: outdata = 32'd9194;
			56343: outdata = 32'd9193;
			56344: outdata = 32'd9192;
			56345: outdata = 32'd9191;
			56346: outdata = 32'd9190;
			56347: outdata = 32'd9189;
			56348: outdata = 32'd9188;
			56349: outdata = 32'd9187;
			56350: outdata = 32'd9186;
			56351: outdata = 32'd9185;
			56352: outdata = 32'd9184;
			56353: outdata = 32'd9183;
			56354: outdata = 32'd9182;
			56355: outdata = 32'd9181;
			56356: outdata = 32'd9180;
			56357: outdata = 32'd9179;
			56358: outdata = 32'd9178;
			56359: outdata = 32'd9177;
			56360: outdata = 32'd9176;
			56361: outdata = 32'd9175;
			56362: outdata = 32'd9174;
			56363: outdata = 32'd9173;
			56364: outdata = 32'd9172;
			56365: outdata = 32'd9171;
			56366: outdata = 32'd9170;
			56367: outdata = 32'd9169;
			56368: outdata = 32'd9168;
			56369: outdata = 32'd9167;
			56370: outdata = 32'd9166;
			56371: outdata = 32'd9165;
			56372: outdata = 32'd9164;
			56373: outdata = 32'd9163;
			56374: outdata = 32'd9162;
			56375: outdata = 32'd9161;
			56376: outdata = 32'd9160;
			56377: outdata = 32'd9159;
			56378: outdata = 32'd9158;
			56379: outdata = 32'd9157;
			56380: outdata = 32'd9156;
			56381: outdata = 32'd9155;
			56382: outdata = 32'd9154;
			56383: outdata = 32'd9153;
			56384: outdata = 32'd9152;
			56385: outdata = 32'd9151;
			56386: outdata = 32'd9150;
			56387: outdata = 32'd9149;
			56388: outdata = 32'd9148;
			56389: outdata = 32'd9147;
			56390: outdata = 32'd9146;
			56391: outdata = 32'd9145;
			56392: outdata = 32'd9144;
			56393: outdata = 32'd9143;
			56394: outdata = 32'd9142;
			56395: outdata = 32'd9141;
			56396: outdata = 32'd9140;
			56397: outdata = 32'd9139;
			56398: outdata = 32'd9138;
			56399: outdata = 32'd9137;
			56400: outdata = 32'd9136;
			56401: outdata = 32'd9135;
			56402: outdata = 32'd9134;
			56403: outdata = 32'd9133;
			56404: outdata = 32'd9132;
			56405: outdata = 32'd9131;
			56406: outdata = 32'd9130;
			56407: outdata = 32'd9129;
			56408: outdata = 32'd9128;
			56409: outdata = 32'd9127;
			56410: outdata = 32'd9126;
			56411: outdata = 32'd9125;
			56412: outdata = 32'd9124;
			56413: outdata = 32'd9123;
			56414: outdata = 32'd9122;
			56415: outdata = 32'd9121;
			56416: outdata = 32'd9120;
			56417: outdata = 32'd9119;
			56418: outdata = 32'd9118;
			56419: outdata = 32'd9117;
			56420: outdata = 32'd9116;
			56421: outdata = 32'd9115;
			56422: outdata = 32'd9114;
			56423: outdata = 32'd9113;
			56424: outdata = 32'd9112;
			56425: outdata = 32'd9111;
			56426: outdata = 32'd9110;
			56427: outdata = 32'd9109;
			56428: outdata = 32'd9108;
			56429: outdata = 32'd9107;
			56430: outdata = 32'd9106;
			56431: outdata = 32'd9105;
			56432: outdata = 32'd9104;
			56433: outdata = 32'd9103;
			56434: outdata = 32'd9102;
			56435: outdata = 32'd9101;
			56436: outdata = 32'd9100;
			56437: outdata = 32'd9099;
			56438: outdata = 32'd9098;
			56439: outdata = 32'd9097;
			56440: outdata = 32'd9096;
			56441: outdata = 32'd9095;
			56442: outdata = 32'd9094;
			56443: outdata = 32'd9093;
			56444: outdata = 32'd9092;
			56445: outdata = 32'd9091;
			56446: outdata = 32'd9090;
			56447: outdata = 32'd9089;
			56448: outdata = 32'd9088;
			56449: outdata = 32'd9087;
			56450: outdata = 32'd9086;
			56451: outdata = 32'd9085;
			56452: outdata = 32'd9084;
			56453: outdata = 32'd9083;
			56454: outdata = 32'd9082;
			56455: outdata = 32'd9081;
			56456: outdata = 32'd9080;
			56457: outdata = 32'd9079;
			56458: outdata = 32'd9078;
			56459: outdata = 32'd9077;
			56460: outdata = 32'd9076;
			56461: outdata = 32'd9075;
			56462: outdata = 32'd9074;
			56463: outdata = 32'd9073;
			56464: outdata = 32'd9072;
			56465: outdata = 32'd9071;
			56466: outdata = 32'd9070;
			56467: outdata = 32'd9069;
			56468: outdata = 32'd9068;
			56469: outdata = 32'd9067;
			56470: outdata = 32'd9066;
			56471: outdata = 32'd9065;
			56472: outdata = 32'd9064;
			56473: outdata = 32'd9063;
			56474: outdata = 32'd9062;
			56475: outdata = 32'd9061;
			56476: outdata = 32'd9060;
			56477: outdata = 32'd9059;
			56478: outdata = 32'd9058;
			56479: outdata = 32'd9057;
			56480: outdata = 32'd9056;
			56481: outdata = 32'd9055;
			56482: outdata = 32'd9054;
			56483: outdata = 32'd9053;
			56484: outdata = 32'd9052;
			56485: outdata = 32'd9051;
			56486: outdata = 32'd9050;
			56487: outdata = 32'd9049;
			56488: outdata = 32'd9048;
			56489: outdata = 32'd9047;
			56490: outdata = 32'd9046;
			56491: outdata = 32'd9045;
			56492: outdata = 32'd9044;
			56493: outdata = 32'd9043;
			56494: outdata = 32'd9042;
			56495: outdata = 32'd9041;
			56496: outdata = 32'd9040;
			56497: outdata = 32'd9039;
			56498: outdata = 32'd9038;
			56499: outdata = 32'd9037;
			56500: outdata = 32'd9036;
			56501: outdata = 32'd9035;
			56502: outdata = 32'd9034;
			56503: outdata = 32'd9033;
			56504: outdata = 32'd9032;
			56505: outdata = 32'd9031;
			56506: outdata = 32'd9030;
			56507: outdata = 32'd9029;
			56508: outdata = 32'd9028;
			56509: outdata = 32'd9027;
			56510: outdata = 32'd9026;
			56511: outdata = 32'd9025;
			56512: outdata = 32'd9024;
			56513: outdata = 32'd9023;
			56514: outdata = 32'd9022;
			56515: outdata = 32'd9021;
			56516: outdata = 32'd9020;
			56517: outdata = 32'd9019;
			56518: outdata = 32'd9018;
			56519: outdata = 32'd9017;
			56520: outdata = 32'd9016;
			56521: outdata = 32'd9015;
			56522: outdata = 32'd9014;
			56523: outdata = 32'd9013;
			56524: outdata = 32'd9012;
			56525: outdata = 32'd9011;
			56526: outdata = 32'd9010;
			56527: outdata = 32'd9009;
			56528: outdata = 32'd9008;
			56529: outdata = 32'd9007;
			56530: outdata = 32'd9006;
			56531: outdata = 32'd9005;
			56532: outdata = 32'd9004;
			56533: outdata = 32'd9003;
			56534: outdata = 32'd9002;
			56535: outdata = 32'd9001;
			56536: outdata = 32'd9000;
			56537: outdata = 32'd8999;
			56538: outdata = 32'd8998;
			56539: outdata = 32'd8997;
			56540: outdata = 32'd8996;
			56541: outdata = 32'd8995;
			56542: outdata = 32'd8994;
			56543: outdata = 32'd8993;
			56544: outdata = 32'd8992;
			56545: outdata = 32'd8991;
			56546: outdata = 32'd8990;
			56547: outdata = 32'd8989;
			56548: outdata = 32'd8988;
			56549: outdata = 32'd8987;
			56550: outdata = 32'd8986;
			56551: outdata = 32'd8985;
			56552: outdata = 32'd8984;
			56553: outdata = 32'd8983;
			56554: outdata = 32'd8982;
			56555: outdata = 32'd8981;
			56556: outdata = 32'd8980;
			56557: outdata = 32'd8979;
			56558: outdata = 32'd8978;
			56559: outdata = 32'd8977;
			56560: outdata = 32'd8976;
			56561: outdata = 32'd8975;
			56562: outdata = 32'd8974;
			56563: outdata = 32'd8973;
			56564: outdata = 32'd8972;
			56565: outdata = 32'd8971;
			56566: outdata = 32'd8970;
			56567: outdata = 32'd8969;
			56568: outdata = 32'd8968;
			56569: outdata = 32'd8967;
			56570: outdata = 32'd8966;
			56571: outdata = 32'd8965;
			56572: outdata = 32'd8964;
			56573: outdata = 32'd8963;
			56574: outdata = 32'd8962;
			56575: outdata = 32'd8961;
			56576: outdata = 32'd8960;
			56577: outdata = 32'd8959;
			56578: outdata = 32'd8958;
			56579: outdata = 32'd8957;
			56580: outdata = 32'd8956;
			56581: outdata = 32'd8955;
			56582: outdata = 32'd8954;
			56583: outdata = 32'd8953;
			56584: outdata = 32'd8952;
			56585: outdata = 32'd8951;
			56586: outdata = 32'd8950;
			56587: outdata = 32'd8949;
			56588: outdata = 32'd8948;
			56589: outdata = 32'd8947;
			56590: outdata = 32'd8946;
			56591: outdata = 32'd8945;
			56592: outdata = 32'd8944;
			56593: outdata = 32'd8943;
			56594: outdata = 32'd8942;
			56595: outdata = 32'd8941;
			56596: outdata = 32'd8940;
			56597: outdata = 32'd8939;
			56598: outdata = 32'd8938;
			56599: outdata = 32'd8937;
			56600: outdata = 32'd8936;
			56601: outdata = 32'd8935;
			56602: outdata = 32'd8934;
			56603: outdata = 32'd8933;
			56604: outdata = 32'd8932;
			56605: outdata = 32'd8931;
			56606: outdata = 32'd8930;
			56607: outdata = 32'd8929;
			56608: outdata = 32'd8928;
			56609: outdata = 32'd8927;
			56610: outdata = 32'd8926;
			56611: outdata = 32'd8925;
			56612: outdata = 32'd8924;
			56613: outdata = 32'd8923;
			56614: outdata = 32'd8922;
			56615: outdata = 32'd8921;
			56616: outdata = 32'd8920;
			56617: outdata = 32'd8919;
			56618: outdata = 32'd8918;
			56619: outdata = 32'd8917;
			56620: outdata = 32'd8916;
			56621: outdata = 32'd8915;
			56622: outdata = 32'd8914;
			56623: outdata = 32'd8913;
			56624: outdata = 32'd8912;
			56625: outdata = 32'd8911;
			56626: outdata = 32'd8910;
			56627: outdata = 32'd8909;
			56628: outdata = 32'd8908;
			56629: outdata = 32'd8907;
			56630: outdata = 32'd8906;
			56631: outdata = 32'd8905;
			56632: outdata = 32'd8904;
			56633: outdata = 32'd8903;
			56634: outdata = 32'd8902;
			56635: outdata = 32'd8901;
			56636: outdata = 32'd8900;
			56637: outdata = 32'd8899;
			56638: outdata = 32'd8898;
			56639: outdata = 32'd8897;
			56640: outdata = 32'd8896;
			56641: outdata = 32'd8895;
			56642: outdata = 32'd8894;
			56643: outdata = 32'd8893;
			56644: outdata = 32'd8892;
			56645: outdata = 32'd8891;
			56646: outdata = 32'd8890;
			56647: outdata = 32'd8889;
			56648: outdata = 32'd8888;
			56649: outdata = 32'd8887;
			56650: outdata = 32'd8886;
			56651: outdata = 32'd8885;
			56652: outdata = 32'd8884;
			56653: outdata = 32'd8883;
			56654: outdata = 32'd8882;
			56655: outdata = 32'd8881;
			56656: outdata = 32'd8880;
			56657: outdata = 32'd8879;
			56658: outdata = 32'd8878;
			56659: outdata = 32'd8877;
			56660: outdata = 32'd8876;
			56661: outdata = 32'd8875;
			56662: outdata = 32'd8874;
			56663: outdata = 32'd8873;
			56664: outdata = 32'd8872;
			56665: outdata = 32'd8871;
			56666: outdata = 32'd8870;
			56667: outdata = 32'd8869;
			56668: outdata = 32'd8868;
			56669: outdata = 32'd8867;
			56670: outdata = 32'd8866;
			56671: outdata = 32'd8865;
			56672: outdata = 32'd8864;
			56673: outdata = 32'd8863;
			56674: outdata = 32'd8862;
			56675: outdata = 32'd8861;
			56676: outdata = 32'd8860;
			56677: outdata = 32'd8859;
			56678: outdata = 32'd8858;
			56679: outdata = 32'd8857;
			56680: outdata = 32'd8856;
			56681: outdata = 32'd8855;
			56682: outdata = 32'd8854;
			56683: outdata = 32'd8853;
			56684: outdata = 32'd8852;
			56685: outdata = 32'd8851;
			56686: outdata = 32'd8850;
			56687: outdata = 32'd8849;
			56688: outdata = 32'd8848;
			56689: outdata = 32'd8847;
			56690: outdata = 32'd8846;
			56691: outdata = 32'd8845;
			56692: outdata = 32'd8844;
			56693: outdata = 32'd8843;
			56694: outdata = 32'd8842;
			56695: outdata = 32'd8841;
			56696: outdata = 32'd8840;
			56697: outdata = 32'd8839;
			56698: outdata = 32'd8838;
			56699: outdata = 32'd8837;
			56700: outdata = 32'd8836;
			56701: outdata = 32'd8835;
			56702: outdata = 32'd8834;
			56703: outdata = 32'd8833;
			56704: outdata = 32'd8832;
			56705: outdata = 32'd8831;
			56706: outdata = 32'd8830;
			56707: outdata = 32'd8829;
			56708: outdata = 32'd8828;
			56709: outdata = 32'd8827;
			56710: outdata = 32'd8826;
			56711: outdata = 32'd8825;
			56712: outdata = 32'd8824;
			56713: outdata = 32'd8823;
			56714: outdata = 32'd8822;
			56715: outdata = 32'd8821;
			56716: outdata = 32'd8820;
			56717: outdata = 32'd8819;
			56718: outdata = 32'd8818;
			56719: outdata = 32'd8817;
			56720: outdata = 32'd8816;
			56721: outdata = 32'd8815;
			56722: outdata = 32'd8814;
			56723: outdata = 32'd8813;
			56724: outdata = 32'd8812;
			56725: outdata = 32'd8811;
			56726: outdata = 32'd8810;
			56727: outdata = 32'd8809;
			56728: outdata = 32'd8808;
			56729: outdata = 32'd8807;
			56730: outdata = 32'd8806;
			56731: outdata = 32'd8805;
			56732: outdata = 32'd8804;
			56733: outdata = 32'd8803;
			56734: outdata = 32'd8802;
			56735: outdata = 32'd8801;
			56736: outdata = 32'd8800;
			56737: outdata = 32'd8799;
			56738: outdata = 32'd8798;
			56739: outdata = 32'd8797;
			56740: outdata = 32'd8796;
			56741: outdata = 32'd8795;
			56742: outdata = 32'd8794;
			56743: outdata = 32'd8793;
			56744: outdata = 32'd8792;
			56745: outdata = 32'd8791;
			56746: outdata = 32'd8790;
			56747: outdata = 32'd8789;
			56748: outdata = 32'd8788;
			56749: outdata = 32'd8787;
			56750: outdata = 32'd8786;
			56751: outdata = 32'd8785;
			56752: outdata = 32'd8784;
			56753: outdata = 32'd8783;
			56754: outdata = 32'd8782;
			56755: outdata = 32'd8781;
			56756: outdata = 32'd8780;
			56757: outdata = 32'd8779;
			56758: outdata = 32'd8778;
			56759: outdata = 32'd8777;
			56760: outdata = 32'd8776;
			56761: outdata = 32'd8775;
			56762: outdata = 32'd8774;
			56763: outdata = 32'd8773;
			56764: outdata = 32'd8772;
			56765: outdata = 32'd8771;
			56766: outdata = 32'd8770;
			56767: outdata = 32'd8769;
			56768: outdata = 32'd8768;
			56769: outdata = 32'd8767;
			56770: outdata = 32'd8766;
			56771: outdata = 32'd8765;
			56772: outdata = 32'd8764;
			56773: outdata = 32'd8763;
			56774: outdata = 32'd8762;
			56775: outdata = 32'd8761;
			56776: outdata = 32'd8760;
			56777: outdata = 32'd8759;
			56778: outdata = 32'd8758;
			56779: outdata = 32'd8757;
			56780: outdata = 32'd8756;
			56781: outdata = 32'd8755;
			56782: outdata = 32'd8754;
			56783: outdata = 32'd8753;
			56784: outdata = 32'd8752;
			56785: outdata = 32'd8751;
			56786: outdata = 32'd8750;
			56787: outdata = 32'd8749;
			56788: outdata = 32'd8748;
			56789: outdata = 32'd8747;
			56790: outdata = 32'd8746;
			56791: outdata = 32'd8745;
			56792: outdata = 32'd8744;
			56793: outdata = 32'd8743;
			56794: outdata = 32'd8742;
			56795: outdata = 32'd8741;
			56796: outdata = 32'd8740;
			56797: outdata = 32'd8739;
			56798: outdata = 32'd8738;
			56799: outdata = 32'd8737;
			56800: outdata = 32'd8736;
			56801: outdata = 32'd8735;
			56802: outdata = 32'd8734;
			56803: outdata = 32'd8733;
			56804: outdata = 32'd8732;
			56805: outdata = 32'd8731;
			56806: outdata = 32'd8730;
			56807: outdata = 32'd8729;
			56808: outdata = 32'd8728;
			56809: outdata = 32'd8727;
			56810: outdata = 32'd8726;
			56811: outdata = 32'd8725;
			56812: outdata = 32'd8724;
			56813: outdata = 32'd8723;
			56814: outdata = 32'd8722;
			56815: outdata = 32'd8721;
			56816: outdata = 32'd8720;
			56817: outdata = 32'd8719;
			56818: outdata = 32'd8718;
			56819: outdata = 32'd8717;
			56820: outdata = 32'd8716;
			56821: outdata = 32'd8715;
			56822: outdata = 32'd8714;
			56823: outdata = 32'd8713;
			56824: outdata = 32'd8712;
			56825: outdata = 32'd8711;
			56826: outdata = 32'd8710;
			56827: outdata = 32'd8709;
			56828: outdata = 32'd8708;
			56829: outdata = 32'd8707;
			56830: outdata = 32'd8706;
			56831: outdata = 32'd8705;
			56832: outdata = 32'd8704;
			56833: outdata = 32'd8703;
			56834: outdata = 32'd8702;
			56835: outdata = 32'd8701;
			56836: outdata = 32'd8700;
			56837: outdata = 32'd8699;
			56838: outdata = 32'd8698;
			56839: outdata = 32'd8697;
			56840: outdata = 32'd8696;
			56841: outdata = 32'd8695;
			56842: outdata = 32'd8694;
			56843: outdata = 32'd8693;
			56844: outdata = 32'd8692;
			56845: outdata = 32'd8691;
			56846: outdata = 32'd8690;
			56847: outdata = 32'd8689;
			56848: outdata = 32'd8688;
			56849: outdata = 32'd8687;
			56850: outdata = 32'd8686;
			56851: outdata = 32'd8685;
			56852: outdata = 32'd8684;
			56853: outdata = 32'd8683;
			56854: outdata = 32'd8682;
			56855: outdata = 32'd8681;
			56856: outdata = 32'd8680;
			56857: outdata = 32'd8679;
			56858: outdata = 32'd8678;
			56859: outdata = 32'd8677;
			56860: outdata = 32'd8676;
			56861: outdata = 32'd8675;
			56862: outdata = 32'd8674;
			56863: outdata = 32'd8673;
			56864: outdata = 32'd8672;
			56865: outdata = 32'd8671;
			56866: outdata = 32'd8670;
			56867: outdata = 32'd8669;
			56868: outdata = 32'd8668;
			56869: outdata = 32'd8667;
			56870: outdata = 32'd8666;
			56871: outdata = 32'd8665;
			56872: outdata = 32'd8664;
			56873: outdata = 32'd8663;
			56874: outdata = 32'd8662;
			56875: outdata = 32'd8661;
			56876: outdata = 32'd8660;
			56877: outdata = 32'd8659;
			56878: outdata = 32'd8658;
			56879: outdata = 32'd8657;
			56880: outdata = 32'd8656;
			56881: outdata = 32'd8655;
			56882: outdata = 32'd8654;
			56883: outdata = 32'd8653;
			56884: outdata = 32'd8652;
			56885: outdata = 32'd8651;
			56886: outdata = 32'd8650;
			56887: outdata = 32'd8649;
			56888: outdata = 32'd8648;
			56889: outdata = 32'd8647;
			56890: outdata = 32'd8646;
			56891: outdata = 32'd8645;
			56892: outdata = 32'd8644;
			56893: outdata = 32'd8643;
			56894: outdata = 32'd8642;
			56895: outdata = 32'd8641;
			56896: outdata = 32'd8640;
			56897: outdata = 32'd8639;
			56898: outdata = 32'd8638;
			56899: outdata = 32'd8637;
			56900: outdata = 32'd8636;
			56901: outdata = 32'd8635;
			56902: outdata = 32'd8634;
			56903: outdata = 32'd8633;
			56904: outdata = 32'd8632;
			56905: outdata = 32'd8631;
			56906: outdata = 32'd8630;
			56907: outdata = 32'd8629;
			56908: outdata = 32'd8628;
			56909: outdata = 32'd8627;
			56910: outdata = 32'd8626;
			56911: outdata = 32'd8625;
			56912: outdata = 32'd8624;
			56913: outdata = 32'd8623;
			56914: outdata = 32'd8622;
			56915: outdata = 32'd8621;
			56916: outdata = 32'd8620;
			56917: outdata = 32'd8619;
			56918: outdata = 32'd8618;
			56919: outdata = 32'd8617;
			56920: outdata = 32'd8616;
			56921: outdata = 32'd8615;
			56922: outdata = 32'd8614;
			56923: outdata = 32'd8613;
			56924: outdata = 32'd8612;
			56925: outdata = 32'd8611;
			56926: outdata = 32'd8610;
			56927: outdata = 32'd8609;
			56928: outdata = 32'd8608;
			56929: outdata = 32'd8607;
			56930: outdata = 32'd8606;
			56931: outdata = 32'd8605;
			56932: outdata = 32'd8604;
			56933: outdata = 32'd8603;
			56934: outdata = 32'd8602;
			56935: outdata = 32'd8601;
			56936: outdata = 32'd8600;
			56937: outdata = 32'd8599;
			56938: outdata = 32'd8598;
			56939: outdata = 32'd8597;
			56940: outdata = 32'd8596;
			56941: outdata = 32'd8595;
			56942: outdata = 32'd8594;
			56943: outdata = 32'd8593;
			56944: outdata = 32'd8592;
			56945: outdata = 32'd8591;
			56946: outdata = 32'd8590;
			56947: outdata = 32'd8589;
			56948: outdata = 32'd8588;
			56949: outdata = 32'd8587;
			56950: outdata = 32'd8586;
			56951: outdata = 32'd8585;
			56952: outdata = 32'd8584;
			56953: outdata = 32'd8583;
			56954: outdata = 32'd8582;
			56955: outdata = 32'd8581;
			56956: outdata = 32'd8580;
			56957: outdata = 32'd8579;
			56958: outdata = 32'd8578;
			56959: outdata = 32'd8577;
			56960: outdata = 32'd8576;
			56961: outdata = 32'd8575;
			56962: outdata = 32'd8574;
			56963: outdata = 32'd8573;
			56964: outdata = 32'd8572;
			56965: outdata = 32'd8571;
			56966: outdata = 32'd8570;
			56967: outdata = 32'd8569;
			56968: outdata = 32'd8568;
			56969: outdata = 32'd8567;
			56970: outdata = 32'd8566;
			56971: outdata = 32'd8565;
			56972: outdata = 32'd8564;
			56973: outdata = 32'd8563;
			56974: outdata = 32'd8562;
			56975: outdata = 32'd8561;
			56976: outdata = 32'd8560;
			56977: outdata = 32'd8559;
			56978: outdata = 32'd8558;
			56979: outdata = 32'd8557;
			56980: outdata = 32'd8556;
			56981: outdata = 32'd8555;
			56982: outdata = 32'd8554;
			56983: outdata = 32'd8553;
			56984: outdata = 32'd8552;
			56985: outdata = 32'd8551;
			56986: outdata = 32'd8550;
			56987: outdata = 32'd8549;
			56988: outdata = 32'd8548;
			56989: outdata = 32'd8547;
			56990: outdata = 32'd8546;
			56991: outdata = 32'd8545;
			56992: outdata = 32'd8544;
			56993: outdata = 32'd8543;
			56994: outdata = 32'd8542;
			56995: outdata = 32'd8541;
			56996: outdata = 32'd8540;
			56997: outdata = 32'd8539;
			56998: outdata = 32'd8538;
			56999: outdata = 32'd8537;
			57000: outdata = 32'd8536;
			57001: outdata = 32'd8535;
			57002: outdata = 32'd8534;
			57003: outdata = 32'd8533;
			57004: outdata = 32'd8532;
			57005: outdata = 32'd8531;
			57006: outdata = 32'd8530;
			57007: outdata = 32'd8529;
			57008: outdata = 32'd8528;
			57009: outdata = 32'd8527;
			57010: outdata = 32'd8526;
			57011: outdata = 32'd8525;
			57012: outdata = 32'd8524;
			57013: outdata = 32'd8523;
			57014: outdata = 32'd8522;
			57015: outdata = 32'd8521;
			57016: outdata = 32'd8520;
			57017: outdata = 32'd8519;
			57018: outdata = 32'd8518;
			57019: outdata = 32'd8517;
			57020: outdata = 32'd8516;
			57021: outdata = 32'd8515;
			57022: outdata = 32'd8514;
			57023: outdata = 32'd8513;
			57024: outdata = 32'd8512;
			57025: outdata = 32'd8511;
			57026: outdata = 32'd8510;
			57027: outdata = 32'd8509;
			57028: outdata = 32'd8508;
			57029: outdata = 32'd8507;
			57030: outdata = 32'd8506;
			57031: outdata = 32'd8505;
			57032: outdata = 32'd8504;
			57033: outdata = 32'd8503;
			57034: outdata = 32'd8502;
			57035: outdata = 32'd8501;
			57036: outdata = 32'd8500;
			57037: outdata = 32'd8499;
			57038: outdata = 32'd8498;
			57039: outdata = 32'd8497;
			57040: outdata = 32'd8496;
			57041: outdata = 32'd8495;
			57042: outdata = 32'd8494;
			57043: outdata = 32'd8493;
			57044: outdata = 32'd8492;
			57045: outdata = 32'd8491;
			57046: outdata = 32'd8490;
			57047: outdata = 32'd8489;
			57048: outdata = 32'd8488;
			57049: outdata = 32'd8487;
			57050: outdata = 32'd8486;
			57051: outdata = 32'd8485;
			57052: outdata = 32'd8484;
			57053: outdata = 32'd8483;
			57054: outdata = 32'd8482;
			57055: outdata = 32'd8481;
			57056: outdata = 32'd8480;
			57057: outdata = 32'd8479;
			57058: outdata = 32'd8478;
			57059: outdata = 32'd8477;
			57060: outdata = 32'd8476;
			57061: outdata = 32'd8475;
			57062: outdata = 32'd8474;
			57063: outdata = 32'd8473;
			57064: outdata = 32'd8472;
			57065: outdata = 32'd8471;
			57066: outdata = 32'd8470;
			57067: outdata = 32'd8469;
			57068: outdata = 32'd8468;
			57069: outdata = 32'd8467;
			57070: outdata = 32'd8466;
			57071: outdata = 32'd8465;
			57072: outdata = 32'd8464;
			57073: outdata = 32'd8463;
			57074: outdata = 32'd8462;
			57075: outdata = 32'd8461;
			57076: outdata = 32'd8460;
			57077: outdata = 32'd8459;
			57078: outdata = 32'd8458;
			57079: outdata = 32'd8457;
			57080: outdata = 32'd8456;
			57081: outdata = 32'd8455;
			57082: outdata = 32'd8454;
			57083: outdata = 32'd8453;
			57084: outdata = 32'd8452;
			57085: outdata = 32'd8451;
			57086: outdata = 32'd8450;
			57087: outdata = 32'd8449;
			57088: outdata = 32'd8448;
			57089: outdata = 32'd8447;
			57090: outdata = 32'd8446;
			57091: outdata = 32'd8445;
			57092: outdata = 32'd8444;
			57093: outdata = 32'd8443;
			57094: outdata = 32'd8442;
			57095: outdata = 32'd8441;
			57096: outdata = 32'd8440;
			57097: outdata = 32'd8439;
			57098: outdata = 32'd8438;
			57099: outdata = 32'd8437;
			57100: outdata = 32'd8436;
			57101: outdata = 32'd8435;
			57102: outdata = 32'd8434;
			57103: outdata = 32'd8433;
			57104: outdata = 32'd8432;
			57105: outdata = 32'd8431;
			57106: outdata = 32'd8430;
			57107: outdata = 32'd8429;
			57108: outdata = 32'd8428;
			57109: outdata = 32'd8427;
			57110: outdata = 32'd8426;
			57111: outdata = 32'd8425;
			57112: outdata = 32'd8424;
			57113: outdata = 32'd8423;
			57114: outdata = 32'd8422;
			57115: outdata = 32'd8421;
			57116: outdata = 32'd8420;
			57117: outdata = 32'd8419;
			57118: outdata = 32'd8418;
			57119: outdata = 32'd8417;
			57120: outdata = 32'd8416;
			57121: outdata = 32'd8415;
			57122: outdata = 32'd8414;
			57123: outdata = 32'd8413;
			57124: outdata = 32'd8412;
			57125: outdata = 32'd8411;
			57126: outdata = 32'd8410;
			57127: outdata = 32'd8409;
			57128: outdata = 32'd8408;
			57129: outdata = 32'd8407;
			57130: outdata = 32'd8406;
			57131: outdata = 32'd8405;
			57132: outdata = 32'd8404;
			57133: outdata = 32'd8403;
			57134: outdata = 32'd8402;
			57135: outdata = 32'd8401;
			57136: outdata = 32'd8400;
			57137: outdata = 32'd8399;
			57138: outdata = 32'd8398;
			57139: outdata = 32'd8397;
			57140: outdata = 32'd8396;
			57141: outdata = 32'd8395;
			57142: outdata = 32'd8394;
			57143: outdata = 32'd8393;
			57144: outdata = 32'd8392;
			57145: outdata = 32'd8391;
			57146: outdata = 32'd8390;
			57147: outdata = 32'd8389;
			57148: outdata = 32'd8388;
			57149: outdata = 32'd8387;
			57150: outdata = 32'd8386;
			57151: outdata = 32'd8385;
			57152: outdata = 32'd8384;
			57153: outdata = 32'd8383;
			57154: outdata = 32'd8382;
			57155: outdata = 32'd8381;
			57156: outdata = 32'd8380;
			57157: outdata = 32'd8379;
			57158: outdata = 32'd8378;
			57159: outdata = 32'd8377;
			57160: outdata = 32'd8376;
			57161: outdata = 32'd8375;
			57162: outdata = 32'd8374;
			57163: outdata = 32'd8373;
			57164: outdata = 32'd8372;
			57165: outdata = 32'd8371;
			57166: outdata = 32'd8370;
			57167: outdata = 32'd8369;
			57168: outdata = 32'd8368;
			57169: outdata = 32'd8367;
			57170: outdata = 32'd8366;
			57171: outdata = 32'd8365;
			57172: outdata = 32'd8364;
			57173: outdata = 32'd8363;
			57174: outdata = 32'd8362;
			57175: outdata = 32'd8361;
			57176: outdata = 32'd8360;
			57177: outdata = 32'd8359;
			57178: outdata = 32'd8358;
			57179: outdata = 32'd8357;
			57180: outdata = 32'd8356;
			57181: outdata = 32'd8355;
			57182: outdata = 32'd8354;
			57183: outdata = 32'd8353;
			57184: outdata = 32'd8352;
			57185: outdata = 32'd8351;
			57186: outdata = 32'd8350;
			57187: outdata = 32'd8349;
			57188: outdata = 32'd8348;
			57189: outdata = 32'd8347;
			57190: outdata = 32'd8346;
			57191: outdata = 32'd8345;
			57192: outdata = 32'd8344;
			57193: outdata = 32'd8343;
			57194: outdata = 32'd8342;
			57195: outdata = 32'd8341;
			57196: outdata = 32'd8340;
			57197: outdata = 32'd8339;
			57198: outdata = 32'd8338;
			57199: outdata = 32'd8337;
			57200: outdata = 32'd8336;
			57201: outdata = 32'd8335;
			57202: outdata = 32'd8334;
			57203: outdata = 32'd8333;
			57204: outdata = 32'd8332;
			57205: outdata = 32'd8331;
			57206: outdata = 32'd8330;
			57207: outdata = 32'd8329;
			57208: outdata = 32'd8328;
			57209: outdata = 32'd8327;
			57210: outdata = 32'd8326;
			57211: outdata = 32'd8325;
			57212: outdata = 32'd8324;
			57213: outdata = 32'd8323;
			57214: outdata = 32'd8322;
			57215: outdata = 32'd8321;
			57216: outdata = 32'd8320;
			57217: outdata = 32'd8319;
			57218: outdata = 32'd8318;
			57219: outdata = 32'd8317;
			57220: outdata = 32'd8316;
			57221: outdata = 32'd8315;
			57222: outdata = 32'd8314;
			57223: outdata = 32'd8313;
			57224: outdata = 32'd8312;
			57225: outdata = 32'd8311;
			57226: outdata = 32'd8310;
			57227: outdata = 32'd8309;
			57228: outdata = 32'd8308;
			57229: outdata = 32'd8307;
			57230: outdata = 32'd8306;
			57231: outdata = 32'd8305;
			57232: outdata = 32'd8304;
			57233: outdata = 32'd8303;
			57234: outdata = 32'd8302;
			57235: outdata = 32'd8301;
			57236: outdata = 32'd8300;
			57237: outdata = 32'd8299;
			57238: outdata = 32'd8298;
			57239: outdata = 32'd8297;
			57240: outdata = 32'd8296;
			57241: outdata = 32'd8295;
			57242: outdata = 32'd8294;
			57243: outdata = 32'd8293;
			57244: outdata = 32'd8292;
			57245: outdata = 32'd8291;
			57246: outdata = 32'd8290;
			57247: outdata = 32'd8289;
			57248: outdata = 32'd8288;
			57249: outdata = 32'd8287;
			57250: outdata = 32'd8286;
			57251: outdata = 32'd8285;
			57252: outdata = 32'd8284;
			57253: outdata = 32'd8283;
			57254: outdata = 32'd8282;
			57255: outdata = 32'd8281;
			57256: outdata = 32'd8280;
			57257: outdata = 32'd8279;
			57258: outdata = 32'd8278;
			57259: outdata = 32'd8277;
			57260: outdata = 32'd8276;
			57261: outdata = 32'd8275;
			57262: outdata = 32'd8274;
			57263: outdata = 32'd8273;
			57264: outdata = 32'd8272;
			57265: outdata = 32'd8271;
			57266: outdata = 32'd8270;
			57267: outdata = 32'd8269;
			57268: outdata = 32'd8268;
			57269: outdata = 32'd8267;
			57270: outdata = 32'd8266;
			57271: outdata = 32'd8265;
			57272: outdata = 32'd8264;
			57273: outdata = 32'd8263;
			57274: outdata = 32'd8262;
			57275: outdata = 32'd8261;
			57276: outdata = 32'd8260;
			57277: outdata = 32'd8259;
			57278: outdata = 32'd8258;
			57279: outdata = 32'd8257;
			57280: outdata = 32'd8256;
			57281: outdata = 32'd8255;
			57282: outdata = 32'd8254;
			57283: outdata = 32'd8253;
			57284: outdata = 32'd8252;
			57285: outdata = 32'd8251;
			57286: outdata = 32'd8250;
			57287: outdata = 32'd8249;
			57288: outdata = 32'd8248;
			57289: outdata = 32'd8247;
			57290: outdata = 32'd8246;
			57291: outdata = 32'd8245;
			57292: outdata = 32'd8244;
			57293: outdata = 32'd8243;
			57294: outdata = 32'd8242;
			57295: outdata = 32'd8241;
			57296: outdata = 32'd8240;
			57297: outdata = 32'd8239;
			57298: outdata = 32'd8238;
			57299: outdata = 32'd8237;
			57300: outdata = 32'd8236;
			57301: outdata = 32'd8235;
			57302: outdata = 32'd8234;
			57303: outdata = 32'd8233;
			57304: outdata = 32'd8232;
			57305: outdata = 32'd8231;
			57306: outdata = 32'd8230;
			57307: outdata = 32'd8229;
			57308: outdata = 32'd8228;
			57309: outdata = 32'd8227;
			57310: outdata = 32'd8226;
			57311: outdata = 32'd8225;
			57312: outdata = 32'd8224;
			57313: outdata = 32'd8223;
			57314: outdata = 32'd8222;
			57315: outdata = 32'd8221;
			57316: outdata = 32'd8220;
			57317: outdata = 32'd8219;
			57318: outdata = 32'd8218;
			57319: outdata = 32'd8217;
			57320: outdata = 32'd8216;
			57321: outdata = 32'd8215;
			57322: outdata = 32'd8214;
			57323: outdata = 32'd8213;
			57324: outdata = 32'd8212;
			57325: outdata = 32'd8211;
			57326: outdata = 32'd8210;
			57327: outdata = 32'd8209;
			57328: outdata = 32'd8208;
			57329: outdata = 32'd8207;
			57330: outdata = 32'd8206;
			57331: outdata = 32'd8205;
			57332: outdata = 32'd8204;
			57333: outdata = 32'd8203;
			57334: outdata = 32'd8202;
			57335: outdata = 32'd8201;
			57336: outdata = 32'd8200;
			57337: outdata = 32'd8199;
			57338: outdata = 32'd8198;
			57339: outdata = 32'd8197;
			57340: outdata = 32'd8196;
			57341: outdata = 32'd8195;
			57342: outdata = 32'd8194;
			57343: outdata = 32'd8193;
			57344: outdata = 32'd8192;
			57345: outdata = 32'd8191;
			57346: outdata = 32'd8190;
			57347: outdata = 32'd8189;
			57348: outdata = 32'd8188;
			57349: outdata = 32'd8187;
			57350: outdata = 32'd8186;
			57351: outdata = 32'd8185;
			57352: outdata = 32'd8184;
			57353: outdata = 32'd8183;
			57354: outdata = 32'd8182;
			57355: outdata = 32'd8181;
			57356: outdata = 32'd8180;
			57357: outdata = 32'd8179;
			57358: outdata = 32'd8178;
			57359: outdata = 32'd8177;
			57360: outdata = 32'd8176;
			57361: outdata = 32'd8175;
			57362: outdata = 32'd8174;
			57363: outdata = 32'd8173;
			57364: outdata = 32'd8172;
			57365: outdata = 32'd8171;
			57366: outdata = 32'd8170;
			57367: outdata = 32'd8169;
			57368: outdata = 32'd8168;
			57369: outdata = 32'd8167;
			57370: outdata = 32'd8166;
			57371: outdata = 32'd8165;
			57372: outdata = 32'd8164;
			57373: outdata = 32'd8163;
			57374: outdata = 32'd8162;
			57375: outdata = 32'd8161;
			57376: outdata = 32'd8160;
			57377: outdata = 32'd8159;
			57378: outdata = 32'd8158;
			57379: outdata = 32'd8157;
			57380: outdata = 32'd8156;
			57381: outdata = 32'd8155;
			57382: outdata = 32'd8154;
			57383: outdata = 32'd8153;
			57384: outdata = 32'd8152;
			57385: outdata = 32'd8151;
			57386: outdata = 32'd8150;
			57387: outdata = 32'd8149;
			57388: outdata = 32'd8148;
			57389: outdata = 32'd8147;
			57390: outdata = 32'd8146;
			57391: outdata = 32'd8145;
			57392: outdata = 32'd8144;
			57393: outdata = 32'd8143;
			57394: outdata = 32'd8142;
			57395: outdata = 32'd8141;
			57396: outdata = 32'd8140;
			57397: outdata = 32'd8139;
			57398: outdata = 32'd8138;
			57399: outdata = 32'd8137;
			57400: outdata = 32'd8136;
			57401: outdata = 32'd8135;
			57402: outdata = 32'd8134;
			57403: outdata = 32'd8133;
			57404: outdata = 32'd8132;
			57405: outdata = 32'd8131;
			57406: outdata = 32'd8130;
			57407: outdata = 32'd8129;
			57408: outdata = 32'd8128;
			57409: outdata = 32'd8127;
			57410: outdata = 32'd8126;
			57411: outdata = 32'd8125;
			57412: outdata = 32'd8124;
			57413: outdata = 32'd8123;
			57414: outdata = 32'd8122;
			57415: outdata = 32'd8121;
			57416: outdata = 32'd8120;
			57417: outdata = 32'd8119;
			57418: outdata = 32'd8118;
			57419: outdata = 32'd8117;
			57420: outdata = 32'd8116;
			57421: outdata = 32'd8115;
			57422: outdata = 32'd8114;
			57423: outdata = 32'd8113;
			57424: outdata = 32'd8112;
			57425: outdata = 32'd8111;
			57426: outdata = 32'd8110;
			57427: outdata = 32'd8109;
			57428: outdata = 32'd8108;
			57429: outdata = 32'd8107;
			57430: outdata = 32'd8106;
			57431: outdata = 32'd8105;
			57432: outdata = 32'd8104;
			57433: outdata = 32'd8103;
			57434: outdata = 32'd8102;
			57435: outdata = 32'd8101;
			57436: outdata = 32'd8100;
			57437: outdata = 32'd8099;
			57438: outdata = 32'd8098;
			57439: outdata = 32'd8097;
			57440: outdata = 32'd8096;
			57441: outdata = 32'd8095;
			57442: outdata = 32'd8094;
			57443: outdata = 32'd8093;
			57444: outdata = 32'd8092;
			57445: outdata = 32'd8091;
			57446: outdata = 32'd8090;
			57447: outdata = 32'd8089;
			57448: outdata = 32'd8088;
			57449: outdata = 32'd8087;
			57450: outdata = 32'd8086;
			57451: outdata = 32'd8085;
			57452: outdata = 32'd8084;
			57453: outdata = 32'd8083;
			57454: outdata = 32'd8082;
			57455: outdata = 32'd8081;
			57456: outdata = 32'd8080;
			57457: outdata = 32'd8079;
			57458: outdata = 32'd8078;
			57459: outdata = 32'd8077;
			57460: outdata = 32'd8076;
			57461: outdata = 32'd8075;
			57462: outdata = 32'd8074;
			57463: outdata = 32'd8073;
			57464: outdata = 32'd8072;
			57465: outdata = 32'd8071;
			57466: outdata = 32'd8070;
			57467: outdata = 32'd8069;
			57468: outdata = 32'd8068;
			57469: outdata = 32'd8067;
			57470: outdata = 32'd8066;
			57471: outdata = 32'd8065;
			57472: outdata = 32'd8064;
			57473: outdata = 32'd8063;
			57474: outdata = 32'd8062;
			57475: outdata = 32'd8061;
			57476: outdata = 32'd8060;
			57477: outdata = 32'd8059;
			57478: outdata = 32'd8058;
			57479: outdata = 32'd8057;
			57480: outdata = 32'd8056;
			57481: outdata = 32'd8055;
			57482: outdata = 32'd8054;
			57483: outdata = 32'd8053;
			57484: outdata = 32'd8052;
			57485: outdata = 32'd8051;
			57486: outdata = 32'd8050;
			57487: outdata = 32'd8049;
			57488: outdata = 32'd8048;
			57489: outdata = 32'd8047;
			57490: outdata = 32'd8046;
			57491: outdata = 32'd8045;
			57492: outdata = 32'd8044;
			57493: outdata = 32'd8043;
			57494: outdata = 32'd8042;
			57495: outdata = 32'd8041;
			57496: outdata = 32'd8040;
			57497: outdata = 32'd8039;
			57498: outdata = 32'd8038;
			57499: outdata = 32'd8037;
			57500: outdata = 32'd8036;
			57501: outdata = 32'd8035;
			57502: outdata = 32'd8034;
			57503: outdata = 32'd8033;
			57504: outdata = 32'd8032;
			57505: outdata = 32'd8031;
			57506: outdata = 32'd8030;
			57507: outdata = 32'd8029;
			57508: outdata = 32'd8028;
			57509: outdata = 32'd8027;
			57510: outdata = 32'd8026;
			57511: outdata = 32'd8025;
			57512: outdata = 32'd8024;
			57513: outdata = 32'd8023;
			57514: outdata = 32'd8022;
			57515: outdata = 32'd8021;
			57516: outdata = 32'd8020;
			57517: outdata = 32'd8019;
			57518: outdata = 32'd8018;
			57519: outdata = 32'd8017;
			57520: outdata = 32'd8016;
			57521: outdata = 32'd8015;
			57522: outdata = 32'd8014;
			57523: outdata = 32'd8013;
			57524: outdata = 32'd8012;
			57525: outdata = 32'd8011;
			57526: outdata = 32'd8010;
			57527: outdata = 32'd8009;
			57528: outdata = 32'd8008;
			57529: outdata = 32'd8007;
			57530: outdata = 32'd8006;
			57531: outdata = 32'd8005;
			57532: outdata = 32'd8004;
			57533: outdata = 32'd8003;
			57534: outdata = 32'd8002;
			57535: outdata = 32'd8001;
			57536: outdata = 32'd8000;
			57537: outdata = 32'd7999;
			57538: outdata = 32'd7998;
			57539: outdata = 32'd7997;
			57540: outdata = 32'd7996;
			57541: outdata = 32'd7995;
			57542: outdata = 32'd7994;
			57543: outdata = 32'd7993;
			57544: outdata = 32'd7992;
			57545: outdata = 32'd7991;
			57546: outdata = 32'd7990;
			57547: outdata = 32'd7989;
			57548: outdata = 32'd7988;
			57549: outdata = 32'd7987;
			57550: outdata = 32'd7986;
			57551: outdata = 32'd7985;
			57552: outdata = 32'd7984;
			57553: outdata = 32'd7983;
			57554: outdata = 32'd7982;
			57555: outdata = 32'd7981;
			57556: outdata = 32'd7980;
			57557: outdata = 32'd7979;
			57558: outdata = 32'd7978;
			57559: outdata = 32'd7977;
			57560: outdata = 32'd7976;
			57561: outdata = 32'd7975;
			57562: outdata = 32'd7974;
			57563: outdata = 32'd7973;
			57564: outdata = 32'd7972;
			57565: outdata = 32'd7971;
			57566: outdata = 32'd7970;
			57567: outdata = 32'd7969;
			57568: outdata = 32'd7968;
			57569: outdata = 32'd7967;
			57570: outdata = 32'd7966;
			57571: outdata = 32'd7965;
			57572: outdata = 32'd7964;
			57573: outdata = 32'd7963;
			57574: outdata = 32'd7962;
			57575: outdata = 32'd7961;
			57576: outdata = 32'd7960;
			57577: outdata = 32'd7959;
			57578: outdata = 32'd7958;
			57579: outdata = 32'd7957;
			57580: outdata = 32'd7956;
			57581: outdata = 32'd7955;
			57582: outdata = 32'd7954;
			57583: outdata = 32'd7953;
			57584: outdata = 32'd7952;
			57585: outdata = 32'd7951;
			57586: outdata = 32'd7950;
			57587: outdata = 32'd7949;
			57588: outdata = 32'd7948;
			57589: outdata = 32'd7947;
			57590: outdata = 32'd7946;
			57591: outdata = 32'd7945;
			57592: outdata = 32'd7944;
			57593: outdata = 32'd7943;
			57594: outdata = 32'd7942;
			57595: outdata = 32'd7941;
			57596: outdata = 32'd7940;
			57597: outdata = 32'd7939;
			57598: outdata = 32'd7938;
			57599: outdata = 32'd7937;
			57600: outdata = 32'd7936;
			57601: outdata = 32'd7935;
			57602: outdata = 32'd7934;
			57603: outdata = 32'd7933;
			57604: outdata = 32'd7932;
			57605: outdata = 32'd7931;
			57606: outdata = 32'd7930;
			57607: outdata = 32'd7929;
			57608: outdata = 32'd7928;
			57609: outdata = 32'd7927;
			57610: outdata = 32'd7926;
			57611: outdata = 32'd7925;
			57612: outdata = 32'd7924;
			57613: outdata = 32'd7923;
			57614: outdata = 32'd7922;
			57615: outdata = 32'd7921;
			57616: outdata = 32'd7920;
			57617: outdata = 32'd7919;
			57618: outdata = 32'd7918;
			57619: outdata = 32'd7917;
			57620: outdata = 32'd7916;
			57621: outdata = 32'd7915;
			57622: outdata = 32'd7914;
			57623: outdata = 32'd7913;
			57624: outdata = 32'd7912;
			57625: outdata = 32'd7911;
			57626: outdata = 32'd7910;
			57627: outdata = 32'd7909;
			57628: outdata = 32'd7908;
			57629: outdata = 32'd7907;
			57630: outdata = 32'd7906;
			57631: outdata = 32'd7905;
			57632: outdata = 32'd7904;
			57633: outdata = 32'd7903;
			57634: outdata = 32'd7902;
			57635: outdata = 32'd7901;
			57636: outdata = 32'd7900;
			57637: outdata = 32'd7899;
			57638: outdata = 32'd7898;
			57639: outdata = 32'd7897;
			57640: outdata = 32'd7896;
			57641: outdata = 32'd7895;
			57642: outdata = 32'd7894;
			57643: outdata = 32'd7893;
			57644: outdata = 32'd7892;
			57645: outdata = 32'd7891;
			57646: outdata = 32'd7890;
			57647: outdata = 32'd7889;
			57648: outdata = 32'd7888;
			57649: outdata = 32'd7887;
			57650: outdata = 32'd7886;
			57651: outdata = 32'd7885;
			57652: outdata = 32'd7884;
			57653: outdata = 32'd7883;
			57654: outdata = 32'd7882;
			57655: outdata = 32'd7881;
			57656: outdata = 32'd7880;
			57657: outdata = 32'd7879;
			57658: outdata = 32'd7878;
			57659: outdata = 32'd7877;
			57660: outdata = 32'd7876;
			57661: outdata = 32'd7875;
			57662: outdata = 32'd7874;
			57663: outdata = 32'd7873;
			57664: outdata = 32'd7872;
			57665: outdata = 32'd7871;
			57666: outdata = 32'd7870;
			57667: outdata = 32'd7869;
			57668: outdata = 32'd7868;
			57669: outdata = 32'd7867;
			57670: outdata = 32'd7866;
			57671: outdata = 32'd7865;
			57672: outdata = 32'd7864;
			57673: outdata = 32'd7863;
			57674: outdata = 32'd7862;
			57675: outdata = 32'd7861;
			57676: outdata = 32'd7860;
			57677: outdata = 32'd7859;
			57678: outdata = 32'd7858;
			57679: outdata = 32'd7857;
			57680: outdata = 32'd7856;
			57681: outdata = 32'd7855;
			57682: outdata = 32'd7854;
			57683: outdata = 32'd7853;
			57684: outdata = 32'd7852;
			57685: outdata = 32'd7851;
			57686: outdata = 32'd7850;
			57687: outdata = 32'd7849;
			57688: outdata = 32'd7848;
			57689: outdata = 32'd7847;
			57690: outdata = 32'd7846;
			57691: outdata = 32'd7845;
			57692: outdata = 32'd7844;
			57693: outdata = 32'd7843;
			57694: outdata = 32'd7842;
			57695: outdata = 32'd7841;
			57696: outdata = 32'd7840;
			57697: outdata = 32'd7839;
			57698: outdata = 32'd7838;
			57699: outdata = 32'd7837;
			57700: outdata = 32'd7836;
			57701: outdata = 32'd7835;
			57702: outdata = 32'd7834;
			57703: outdata = 32'd7833;
			57704: outdata = 32'd7832;
			57705: outdata = 32'd7831;
			57706: outdata = 32'd7830;
			57707: outdata = 32'd7829;
			57708: outdata = 32'd7828;
			57709: outdata = 32'd7827;
			57710: outdata = 32'd7826;
			57711: outdata = 32'd7825;
			57712: outdata = 32'd7824;
			57713: outdata = 32'd7823;
			57714: outdata = 32'd7822;
			57715: outdata = 32'd7821;
			57716: outdata = 32'd7820;
			57717: outdata = 32'd7819;
			57718: outdata = 32'd7818;
			57719: outdata = 32'd7817;
			57720: outdata = 32'd7816;
			57721: outdata = 32'd7815;
			57722: outdata = 32'd7814;
			57723: outdata = 32'd7813;
			57724: outdata = 32'd7812;
			57725: outdata = 32'd7811;
			57726: outdata = 32'd7810;
			57727: outdata = 32'd7809;
			57728: outdata = 32'd7808;
			57729: outdata = 32'd7807;
			57730: outdata = 32'd7806;
			57731: outdata = 32'd7805;
			57732: outdata = 32'd7804;
			57733: outdata = 32'd7803;
			57734: outdata = 32'd7802;
			57735: outdata = 32'd7801;
			57736: outdata = 32'd7800;
			57737: outdata = 32'd7799;
			57738: outdata = 32'd7798;
			57739: outdata = 32'd7797;
			57740: outdata = 32'd7796;
			57741: outdata = 32'd7795;
			57742: outdata = 32'd7794;
			57743: outdata = 32'd7793;
			57744: outdata = 32'd7792;
			57745: outdata = 32'd7791;
			57746: outdata = 32'd7790;
			57747: outdata = 32'd7789;
			57748: outdata = 32'd7788;
			57749: outdata = 32'd7787;
			57750: outdata = 32'd7786;
			57751: outdata = 32'd7785;
			57752: outdata = 32'd7784;
			57753: outdata = 32'd7783;
			57754: outdata = 32'd7782;
			57755: outdata = 32'd7781;
			57756: outdata = 32'd7780;
			57757: outdata = 32'd7779;
			57758: outdata = 32'd7778;
			57759: outdata = 32'd7777;
			57760: outdata = 32'd7776;
			57761: outdata = 32'd7775;
			57762: outdata = 32'd7774;
			57763: outdata = 32'd7773;
			57764: outdata = 32'd7772;
			57765: outdata = 32'd7771;
			57766: outdata = 32'd7770;
			57767: outdata = 32'd7769;
			57768: outdata = 32'd7768;
			57769: outdata = 32'd7767;
			57770: outdata = 32'd7766;
			57771: outdata = 32'd7765;
			57772: outdata = 32'd7764;
			57773: outdata = 32'd7763;
			57774: outdata = 32'd7762;
			57775: outdata = 32'd7761;
			57776: outdata = 32'd7760;
			57777: outdata = 32'd7759;
			57778: outdata = 32'd7758;
			57779: outdata = 32'd7757;
			57780: outdata = 32'd7756;
			57781: outdata = 32'd7755;
			57782: outdata = 32'd7754;
			57783: outdata = 32'd7753;
			57784: outdata = 32'd7752;
			57785: outdata = 32'd7751;
			57786: outdata = 32'd7750;
			57787: outdata = 32'd7749;
			57788: outdata = 32'd7748;
			57789: outdata = 32'd7747;
			57790: outdata = 32'd7746;
			57791: outdata = 32'd7745;
			57792: outdata = 32'd7744;
			57793: outdata = 32'd7743;
			57794: outdata = 32'd7742;
			57795: outdata = 32'd7741;
			57796: outdata = 32'd7740;
			57797: outdata = 32'd7739;
			57798: outdata = 32'd7738;
			57799: outdata = 32'd7737;
			57800: outdata = 32'd7736;
			57801: outdata = 32'd7735;
			57802: outdata = 32'd7734;
			57803: outdata = 32'd7733;
			57804: outdata = 32'd7732;
			57805: outdata = 32'd7731;
			57806: outdata = 32'd7730;
			57807: outdata = 32'd7729;
			57808: outdata = 32'd7728;
			57809: outdata = 32'd7727;
			57810: outdata = 32'd7726;
			57811: outdata = 32'd7725;
			57812: outdata = 32'd7724;
			57813: outdata = 32'd7723;
			57814: outdata = 32'd7722;
			57815: outdata = 32'd7721;
			57816: outdata = 32'd7720;
			57817: outdata = 32'd7719;
			57818: outdata = 32'd7718;
			57819: outdata = 32'd7717;
			57820: outdata = 32'd7716;
			57821: outdata = 32'd7715;
			57822: outdata = 32'd7714;
			57823: outdata = 32'd7713;
			57824: outdata = 32'd7712;
			57825: outdata = 32'd7711;
			57826: outdata = 32'd7710;
			57827: outdata = 32'd7709;
			57828: outdata = 32'd7708;
			57829: outdata = 32'd7707;
			57830: outdata = 32'd7706;
			57831: outdata = 32'd7705;
			57832: outdata = 32'd7704;
			57833: outdata = 32'd7703;
			57834: outdata = 32'd7702;
			57835: outdata = 32'd7701;
			57836: outdata = 32'd7700;
			57837: outdata = 32'd7699;
			57838: outdata = 32'd7698;
			57839: outdata = 32'd7697;
			57840: outdata = 32'd7696;
			57841: outdata = 32'd7695;
			57842: outdata = 32'd7694;
			57843: outdata = 32'd7693;
			57844: outdata = 32'd7692;
			57845: outdata = 32'd7691;
			57846: outdata = 32'd7690;
			57847: outdata = 32'd7689;
			57848: outdata = 32'd7688;
			57849: outdata = 32'd7687;
			57850: outdata = 32'd7686;
			57851: outdata = 32'd7685;
			57852: outdata = 32'd7684;
			57853: outdata = 32'd7683;
			57854: outdata = 32'd7682;
			57855: outdata = 32'd7681;
			57856: outdata = 32'd7680;
			57857: outdata = 32'd7679;
			57858: outdata = 32'd7678;
			57859: outdata = 32'd7677;
			57860: outdata = 32'd7676;
			57861: outdata = 32'd7675;
			57862: outdata = 32'd7674;
			57863: outdata = 32'd7673;
			57864: outdata = 32'd7672;
			57865: outdata = 32'd7671;
			57866: outdata = 32'd7670;
			57867: outdata = 32'd7669;
			57868: outdata = 32'd7668;
			57869: outdata = 32'd7667;
			57870: outdata = 32'd7666;
			57871: outdata = 32'd7665;
			57872: outdata = 32'd7664;
			57873: outdata = 32'd7663;
			57874: outdata = 32'd7662;
			57875: outdata = 32'd7661;
			57876: outdata = 32'd7660;
			57877: outdata = 32'd7659;
			57878: outdata = 32'd7658;
			57879: outdata = 32'd7657;
			57880: outdata = 32'd7656;
			57881: outdata = 32'd7655;
			57882: outdata = 32'd7654;
			57883: outdata = 32'd7653;
			57884: outdata = 32'd7652;
			57885: outdata = 32'd7651;
			57886: outdata = 32'd7650;
			57887: outdata = 32'd7649;
			57888: outdata = 32'd7648;
			57889: outdata = 32'd7647;
			57890: outdata = 32'd7646;
			57891: outdata = 32'd7645;
			57892: outdata = 32'd7644;
			57893: outdata = 32'd7643;
			57894: outdata = 32'd7642;
			57895: outdata = 32'd7641;
			57896: outdata = 32'd7640;
			57897: outdata = 32'd7639;
			57898: outdata = 32'd7638;
			57899: outdata = 32'd7637;
			57900: outdata = 32'd7636;
			57901: outdata = 32'd7635;
			57902: outdata = 32'd7634;
			57903: outdata = 32'd7633;
			57904: outdata = 32'd7632;
			57905: outdata = 32'd7631;
			57906: outdata = 32'd7630;
			57907: outdata = 32'd7629;
			57908: outdata = 32'd7628;
			57909: outdata = 32'd7627;
			57910: outdata = 32'd7626;
			57911: outdata = 32'd7625;
			57912: outdata = 32'd7624;
			57913: outdata = 32'd7623;
			57914: outdata = 32'd7622;
			57915: outdata = 32'd7621;
			57916: outdata = 32'd7620;
			57917: outdata = 32'd7619;
			57918: outdata = 32'd7618;
			57919: outdata = 32'd7617;
			57920: outdata = 32'd7616;
			57921: outdata = 32'd7615;
			57922: outdata = 32'd7614;
			57923: outdata = 32'd7613;
			57924: outdata = 32'd7612;
			57925: outdata = 32'd7611;
			57926: outdata = 32'd7610;
			57927: outdata = 32'd7609;
			57928: outdata = 32'd7608;
			57929: outdata = 32'd7607;
			57930: outdata = 32'd7606;
			57931: outdata = 32'd7605;
			57932: outdata = 32'd7604;
			57933: outdata = 32'd7603;
			57934: outdata = 32'd7602;
			57935: outdata = 32'd7601;
			57936: outdata = 32'd7600;
			57937: outdata = 32'd7599;
			57938: outdata = 32'd7598;
			57939: outdata = 32'd7597;
			57940: outdata = 32'd7596;
			57941: outdata = 32'd7595;
			57942: outdata = 32'd7594;
			57943: outdata = 32'd7593;
			57944: outdata = 32'd7592;
			57945: outdata = 32'd7591;
			57946: outdata = 32'd7590;
			57947: outdata = 32'd7589;
			57948: outdata = 32'd7588;
			57949: outdata = 32'd7587;
			57950: outdata = 32'd7586;
			57951: outdata = 32'd7585;
			57952: outdata = 32'd7584;
			57953: outdata = 32'd7583;
			57954: outdata = 32'd7582;
			57955: outdata = 32'd7581;
			57956: outdata = 32'd7580;
			57957: outdata = 32'd7579;
			57958: outdata = 32'd7578;
			57959: outdata = 32'd7577;
			57960: outdata = 32'd7576;
			57961: outdata = 32'd7575;
			57962: outdata = 32'd7574;
			57963: outdata = 32'd7573;
			57964: outdata = 32'd7572;
			57965: outdata = 32'd7571;
			57966: outdata = 32'd7570;
			57967: outdata = 32'd7569;
			57968: outdata = 32'd7568;
			57969: outdata = 32'd7567;
			57970: outdata = 32'd7566;
			57971: outdata = 32'd7565;
			57972: outdata = 32'd7564;
			57973: outdata = 32'd7563;
			57974: outdata = 32'd7562;
			57975: outdata = 32'd7561;
			57976: outdata = 32'd7560;
			57977: outdata = 32'd7559;
			57978: outdata = 32'd7558;
			57979: outdata = 32'd7557;
			57980: outdata = 32'd7556;
			57981: outdata = 32'd7555;
			57982: outdata = 32'd7554;
			57983: outdata = 32'd7553;
			57984: outdata = 32'd7552;
			57985: outdata = 32'd7551;
			57986: outdata = 32'd7550;
			57987: outdata = 32'd7549;
			57988: outdata = 32'd7548;
			57989: outdata = 32'd7547;
			57990: outdata = 32'd7546;
			57991: outdata = 32'd7545;
			57992: outdata = 32'd7544;
			57993: outdata = 32'd7543;
			57994: outdata = 32'd7542;
			57995: outdata = 32'd7541;
			57996: outdata = 32'd7540;
			57997: outdata = 32'd7539;
			57998: outdata = 32'd7538;
			57999: outdata = 32'd7537;
			58000: outdata = 32'd7536;
			58001: outdata = 32'd7535;
			58002: outdata = 32'd7534;
			58003: outdata = 32'd7533;
			58004: outdata = 32'd7532;
			58005: outdata = 32'd7531;
			58006: outdata = 32'd7530;
			58007: outdata = 32'd7529;
			58008: outdata = 32'd7528;
			58009: outdata = 32'd7527;
			58010: outdata = 32'd7526;
			58011: outdata = 32'd7525;
			58012: outdata = 32'd7524;
			58013: outdata = 32'd7523;
			58014: outdata = 32'd7522;
			58015: outdata = 32'd7521;
			58016: outdata = 32'd7520;
			58017: outdata = 32'd7519;
			58018: outdata = 32'd7518;
			58019: outdata = 32'd7517;
			58020: outdata = 32'd7516;
			58021: outdata = 32'd7515;
			58022: outdata = 32'd7514;
			58023: outdata = 32'd7513;
			58024: outdata = 32'd7512;
			58025: outdata = 32'd7511;
			58026: outdata = 32'd7510;
			58027: outdata = 32'd7509;
			58028: outdata = 32'd7508;
			58029: outdata = 32'd7507;
			58030: outdata = 32'd7506;
			58031: outdata = 32'd7505;
			58032: outdata = 32'd7504;
			58033: outdata = 32'd7503;
			58034: outdata = 32'd7502;
			58035: outdata = 32'd7501;
			58036: outdata = 32'd7500;
			58037: outdata = 32'd7499;
			58038: outdata = 32'd7498;
			58039: outdata = 32'd7497;
			58040: outdata = 32'd7496;
			58041: outdata = 32'd7495;
			58042: outdata = 32'd7494;
			58043: outdata = 32'd7493;
			58044: outdata = 32'd7492;
			58045: outdata = 32'd7491;
			58046: outdata = 32'd7490;
			58047: outdata = 32'd7489;
			58048: outdata = 32'd7488;
			58049: outdata = 32'd7487;
			58050: outdata = 32'd7486;
			58051: outdata = 32'd7485;
			58052: outdata = 32'd7484;
			58053: outdata = 32'd7483;
			58054: outdata = 32'd7482;
			58055: outdata = 32'd7481;
			58056: outdata = 32'd7480;
			58057: outdata = 32'd7479;
			58058: outdata = 32'd7478;
			58059: outdata = 32'd7477;
			58060: outdata = 32'd7476;
			58061: outdata = 32'd7475;
			58062: outdata = 32'd7474;
			58063: outdata = 32'd7473;
			58064: outdata = 32'd7472;
			58065: outdata = 32'd7471;
			58066: outdata = 32'd7470;
			58067: outdata = 32'd7469;
			58068: outdata = 32'd7468;
			58069: outdata = 32'd7467;
			58070: outdata = 32'd7466;
			58071: outdata = 32'd7465;
			58072: outdata = 32'd7464;
			58073: outdata = 32'd7463;
			58074: outdata = 32'd7462;
			58075: outdata = 32'd7461;
			58076: outdata = 32'd7460;
			58077: outdata = 32'd7459;
			58078: outdata = 32'd7458;
			58079: outdata = 32'd7457;
			58080: outdata = 32'd7456;
			58081: outdata = 32'd7455;
			58082: outdata = 32'd7454;
			58083: outdata = 32'd7453;
			58084: outdata = 32'd7452;
			58085: outdata = 32'd7451;
			58086: outdata = 32'd7450;
			58087: outdata = 32'd7449;
			58088: outdata = 32'd7448;
			58089: outdata = 32'd7447;
			58090: outdata = 32'd7446;
			58091: outdata = 32'd7445;
			58092: outdata = 32'd7444;
			58093: outdata = 32'd7443;
			58094: outdata = 32'd7442;
			58095: outdata = 32'd7441;
			58096: outdata = 32'd7440;
			58097: outdata = 32'd7439;
			58098: outdata = 32'd7438;
			58099: outdata = 32'd7437;
			58100: outdata = 32'd7436;
			58101: outdata = 32'd7435;
			58102: outdata = 32'd7434;
			58103: outdata = 32'd7433;
			58104: outdata = 32'd7432;
			58105: outdata = 32'd7431;
			58106: outdata = 32'd7430;
			58107: outdata = 32'd7429;
			58108: outdata = 32'd7428;
			58109: outdata = 32'd7427;
			58110: outdata = 32'd7426;
			58111: outdata = 32'd7425;
			58112: outdata = 32'd7424;
			58113: outdata = 32'd7423;
			58114: outdata = 32'd7422;
			58115: outdata = 32'd7421;
			58116: outdata = 32'd7420;
			58117: outdata = 32'd7419;
			58118: outdata = 32'd7418;
			58119: outdata = 32'd7417;
			58120: outdata = 32'd7416;
			58121: outdata = 32'd7415;
			58122: outdata = 32'd7414;
			58123: outdata = 32'd7413;
			58124: outdata = 32'd7412;
			58125: outdata = 32'd7411;
			58126: outdata = 32'd7410;
			58127: outdata = 32'd7409;
			58128: outdata = 32'd7408;
			58129: outdata = 32'd7407;
			58130: outdata = 32'd7406;
			58131: outdata = 32'd7405;
			58132: outdata = 32'd7404;
			58133: outdata = 32'd7403;
			58134: outdata = 32'd7402;
			58135: outdata = 32'd7401;
			58136: outdata = 32'd7400;
			58137: outdata = 32'd7399;
			58138: outdata = 32'd7398;
			58139: outdata = 32'd7397;
			58140: outdata = 32'd7396;
			58141: outdata = 32'd7395;
			58142: outdata = 32'd7394;
			58143: outdata = 32'd7393;
			58144: outdata = 32'd7392;
			58145: outdata = 32'd7391;
			58146: outdata = 32'd7390;
			58147: outdata = 32'd7389;
			58148: outdata = 32'd7388;
			58149: outdata = 32'd7387;
			58150: outdata = 32'd7386;
			58151: outdata = 32'd7385;
			58152: outdata = 32'd7384;
			58153: outdata = 32'd7383;
			58154: outdata = 32'd7382;
			58155: outdata = 32'd7381;
			58156: outdata = 32'd7380;
			58157: outdata = 32'd7379;
			58158: outdata = 32'd7378;
			58159: outdata = 32'd7377;
			58160: outdata = 32'd7376;
			58161: outdata = 32'd7375;
			58162: outdata = 32'd7374;
			58163: outdata = 32'd7373;
			58164: outdata = 32'd7372;
			58165: outdata = 32'd7371;
			58166: outdata = 32'd7370;
			58167: outdata = 32'd7369;
			58168: outdata = 32'd7368;
			58169: outdata = 32'd7367;
			58170: outdata = 32'd7366;
			58171: outdata = 32'd7365;
			58172: outdata = 32'd7364;
			58173: outdata = 32'd7363;
			58174: outdata = 32'd7362;
			58175: outdata = 32'd7361;
			58176: outdata = 32'd7360;
			58177: outdata = 32'd7359;
			58178: outdata = 32'd7358;
			58179: outdata = 32'd7357;
			58180: outdata = 32'd7356;
			58181: outdata = 32'd7355;
			58182: outdata = 32'd7354;
			58183: outdata = 32'd7353;
			58184: outdata = 32'd7352;
			58185: outdata = 32'd7351;
			58186: outdata = 32'd7350;
			58187: outdata = 32'd7349;
			58188: outdata = 32'd7348;
			58189: outdata = 32'd7347;
			58190: outdata = 32'd7346;
			58191: outdata = 32'd7345;
			58192: outdata = 32'd7344;
			58193: outdata = 32'd7343;
			58194: outdata = 32'd7342;
			58195: outdata = 32'd7341;
			58196: outdata = 32'd7340;
			58197: outdata = 32'd7339;
			58198: outdata = 32'd7338;
			58199: outdata = 32'd7337;
			58200: outdata = 32'd7336;
			58201: outdata = 32'd7335;
			58202: outdata = 32'd7334;
			58203: outdata = 32'd7333;
			58204: outdata = 32'd7332;
			58205: outdata = 32'd7331;
			58206: outdata = 32'd7330;
			58207: outdata = 32'd7329;
			58208: outdata = 32'd7328;
			58209: outdata = 32'd7327;
			58210: outdata = 32'd7326;
			58211: outdata = 32'd7325;
			58212: outdata = 32'd7324;
			58213: outdata = 32'd7323;
			58214: outdata = 32'd7322;
			58215: outdata = 32'd7321;
			58216: outdata = 32'd7320;
			58217: outdata = 32'd7319;
			58218: outdata = 32'd7318;
			58219: outdata = 32'd7317;
			58220: outdata = 32'd7316;
			58221: outdata = 32'd7315;
			58222: outdata = 32'd7314;
			58223: outdata = 32'd7313;
			58224: outdata = 32'd7312;
			58225: outdata = 32'd7311;
			58226: outdata = 32'd7310;
			58227: outdata = 32'd7309;
			58228: outdata = 32'd7308;
			58229: outdata = 32'd7307;
			58230: outdata = 32'd7306;
			58231: outdata = 32'd7305;
			58232: outdata = 32'd7304;
			58233: outdata = 32'd7303;
			58234: outdata = 32'd7302;
			58235: outdata = 32'd7301;
			58236: outdata = 32'd7300;
			58237: outdata = 32'd7299;
			58238: outdata = 32'd7298;
			58239: outdata = 32'd7297;
			58240: outdata = 32'd7296;
			58241: outdata = 32'd7295;
			58242: outdata = 32'd7294;
			58243: outdata = 32'd7293;
			58244: outdata = 32'd7292;
			58245: outdata = 32'd7291;
			58246: outdata = 32'd7290;
			58247: outdata = 32'd7289;
			58248: outdata = 32'd7288;
			58249: outdata = 32'd7287;
			58250: outdata = 32'd7286;
			58251: outdata = 32'd7285;
			58252: outdata = 32'd7284;
			58253: outdata = 32'd7283;
			58254: outdata = 32'd7282;
			58255: outdata = 32'd7281;
			58256: outdata = 32'd7280;
			58257: outdata = 32'd7279;
			58258: outdata = 32'd7278;
			58259: outdata = 32'd7277;
			58260: outdata = 32'd7276;
			58261: outdata = 32'd7275;
			58262: outdata = 32'd7274;
			58263: outdata = 32'd7273;
			58264: outdata = 32'd7272;
			58265: outdata = 32'd7271;
			58266: outdata = 32'd7270;
			58267: outdata = 32'd7269;
			58268: outdata = 32'd7268;
			58269: outdata = 32'd7267;
			58270: outdata = 32'd7266;
			58271: outdata = 32'd7265;
			58272: outdata = 32'd7264;
			58273: outdata = 32'd7263;
			58274: outdata = 32'd7262;
			58275: outdata = 32'd7261;
			58276: outdata = 32'd7260;
			58277: outdata = 32'd7259;
			58278: outdata = 32'd7258;
			58279: outdata = 32'd7257;
			58280: outdata = 32'd7256;
			58281: outdata = 32'd7255;
			58282: outdata = 32'd7254;
			58283: outdata = 32'd7253;
			58284: outdata = 32'd7252;
			58285: outdata = 32'd7251;
			58286: outdata = 32'd7250;
			58287: outdata = 32'd7249;
			58288: outdata = 32'd7248;
			58289: outdata = 32'd7247;
			58290: outdata = 32'd7246;
			58291: outdata = 32'd7245;
			58292: outdata = 32'd7244;
			58293: outdata = 32'd7243;
			58294: outdata = 32'd7242;
			58295: outdata = 32'd7241;
			58296: outdata = 32'd7240;
			58297: outdata = 32'd7239;
			58298: outdata = 32'd7238;
			58299: outdata = 32'd7237;
			58300: outdata = 32'd7236;
			58301: outdata = 32'd7235;
			58302: outdata = 32'd7234;
			58303: outdata = 32'd7233;
			58304: outdata = 32'd7232;
			58305: outdata = 32'd7231;
			58306: outdata = 32'd7230;
			58307: outdata = 32'd7229;
			58308: outdata = 32'd7228;
			58309: outdata = 32'd7227;
			58310: outdata = 32'd7226;
			58311: outdata = 32'd7225;
			58312: outdata = 32'd7224;
			58313: outdata = 32'd7223;
			58314: outdata = 32'd7222;
			58315: outdata = 32'd7221;
			58316: outdata = 32'd7220;
			58317: outdata = 32'd7219;
			58318: outdata = 32'd7218;
			58319: outdata = 32'd7217;
			58320: outdata = 32'd7216;
			58321: outdata = 32'd7215;
			58322: outdata = 32'd7214;
			58323: outdata = 32'd7213;
			58324: outdata = 32'd7212;
			58325: outdata = 32'd7211;
			58326: outdata = 32'd7210;
			58327: outdata = 32'd7209;
			58328: outdata = 32'd7208;
			58329: outdata = 32'd7207;
			58330: outdata = 32'd7206;
			58331: outdata = 32'd7205;
			58332: outdata = 32'd7204;
			58333: outdata = 32'd7203;
			58334: outdata = 32'd7202;
			58335: outdata = 32'd7201;
			58336: outdata = 32'd7200;
			58337: outdata = 32'd7199;
			58338: outdata = 32'd7198;
			58339: outdata = 32'd7197;
			58340: outdata = 32'd7196;
			58341: outdata = 32'd7195;
			58342: outdata = 32'd7194;
			58343: outdata = 32'd7193;
			58344: outdata = 32'd7192;
			58345: outdata = 32'd7191;
			58346: outdata = 32'd7190;
			58347: outdata = 32'd7189;
			58348: outdata = 32'd7188;
			58349: outdata = 32'd7187;
			58350: outdata = 32'd7186;
			58351: outdata = 32'd7185;
			58352: outdata = 32'd7184;
			58353: outdata = 32'd7183;
			58354: outdata = 32'd7182;
			58355: outdata = 32'd7181;
			58356: outdata = 32'd7180;
			58357: outdata = 32'd7179;
			58358: outdata = 32'd7178;
			58359: outdata = 32'd7177;
			58360: outdata = 32'd7176;
			58361: outdata = 32'd7175;
			58362: outdata = 32'd7174;
			58363: outdata = 32'd7173;
			58364: outdata = 32'd7172;
			58365: outdata = 32'd7171;
			58366: outdata = 32'd7170;
			58367: outdata = 32'd7169;
			58368: outdata = 32'd7168;
			58369: outdata = 32'd7167;
			58370: outdata = 32'd7166;
			58371: outdata = 32'd7165;
			58372: outdata = 32'd7164;
			58373: outdata = 32'd7163;
			58374: outdata = 32'd7162;
			58375: outdata = 32'd7161;
			58376: outdata = 32'd7160;
			58377: outdata = 32'd7159;
			58378: outdata = 32'd7158;
			58379: outdata = 32'd7157;
			58380: outdata = 32'd7156;
			58381: outdata = 32'd7155;
			58382: outdata = 32'd7154;
			58383: outdata = 32'd7153;
			58384: outdata = 32'd7152;
			58385: outdata = 32'd7151;
			58386: outdata = 32'd7150;
			58387: outdata = 32'd7149;
			58388: outdata = 32'd7148;
			58389: outdata = 32'd7147;
			58390: outdata = 32'd7146;
			58391: outdata = 32'd7145;
			58392: outdata = 32'd7144;
			58393: outdata = 32'd7143;
			58394: outdata = 32'd7142;
			58395: outdata = 32'd7141;
			58396: outdata = 32'd7140;
			58397: outdata = 32'd7139;
			58398: outdata = 32'd7138;
			58399: outdata = 32'd7137;
			58400: outdata = 32'd7136;
			58401: outdata = 32'd7135;
			58402: outdata = 32'd7134;
			58403: outdata = 32'd7133;
			58404: outdata = 32'd7132;
			58405: outdata = 32'd7131;
			58406: outdata = 32'd7130;
			58407: outdata = 32'd7129;
			58408: outdata = 32'd7128;
			58409: outdata = 32'd7127;
			58410: outdata = 32'd7126;
			58411: outdata = 32'd7125;
			58412: outdata = 32'd7124;
			58413: outdata = 32'd7123;
			58414: outdata = 32'd7122;
			58415: outdata = 32'd7121;
			58416: outdata = 32'd7120;
			58417: outdata = 32'd7119;
			58418: outdata = 32'd7118;
			58419: outdata = 32'd7117;
			58420: outdata = 32'd7116;
			58421: outdata = 32'd7115;
			58422: outdata = 32'd7114;
			58423: outdata = 32'd7113;
			58424: outdata = 32'd7112;
			58425: outdata = 32'd7111;
			58426: outdata = 32'd7110;
			58427: outdata = 32'd7109;
			58428: outdata = 32'd7108;
			58429: outdata = 32'd7107;
			58430: outdata = 32'd7106;
			58431: outdata = 32'd7105;
			58432: outdata = 32'd7104;
			58433: outdata = 32'd7103;
			58434: outdata = 32'd7102;
			58435: outdata = 32'd7101;
			58436: outdata = 32'd7100;
			58437: outdata = 32'd7099;
			58438: outdata = 32'd7098;
			58439: outdata = 32'd7097;
			58440: outdata = 32'd7096;
			58441: outdata = 32'd7095;
			58442: outdata = 32'd7094;
			58443: outdata = 32'd7093;
			58444: outdata = 32'd7092;
			58445: outdata = 32'd7091;
			58446: outdata = 32'd7090;
			58447: outdata = 32'd7089;
			58448: outdata = 32'd7088;
			58449: outdata = 32'd7087;
			58450: outdata = 32'd7086;
			58451: outdata = 32'd7085;
			58452: outdata = 32'd7084;
			58453: outdata = 32'd7083;
			58454: outdata = 32'd7082;
			58455: outdata = 32'd7081;
			58456: outdata = 32'd7080;
			58457: outdata = 32'd7079;
			58458: outdata = 32'd7078;
			58459: outdata = 32'd7077;
			58460: outdata = 32'd7076;
			58461: outdata = 32'd7075;
			58462: outdata = 32'd7074;
			58463: outdata = 32'd7073;
			58464: outdata = 32'd7072;
			58465: outdata = 32'd7071;
			58466: outdata = 32'd7070;
			58467: outdata = 32'd7069;
			58468: outdata = 32'd7068;
			58469: outdata = 32'd7067;
			58470: outdata = 32'd7066;
			58471: outdata = 32'd7065;
			58472: outdata = 32'd7064;
			58473: outdata = 32'd7063;
			58474: outdata = 32'd7062;
			58475: outdata = 32'd7061;
			58476: outdata = 32'd7060;
			58477: outdata = 32'd7059;
			58478: outdata = 32'd7058;
			58479: outdata = 32'd7057;
			58480: outdata = 32'd7056;
			58481: outdata = 32'd7055;
			58482: outdata = 32'd7054;
			58483: outdata = 32'd7053;
			58484: outdata = 32'd7052;
			58485: outdata = 32'd7051;
			58486: outdata = 32'd7050;
			58487: outdata = 32'd7049;
			58488: outdata = 32'd7048;
			58489: outdata = 32'd7047;
			58490: outdata = 32'd7046;
			58491: outdata = 32'd7045;
			58492: outdata = 32'd7044;
			58493: outdata = 32'd7043;
			58494: outdata = 32'd7042;
			58495: outdata = 32'd7041;
			58496: outdata = 32'd7040;
			58497: outdata = 32'd7039;
			58498: outdata = 32'd7038;
			58499: outdata = 32'd7037;
			58500: outdata = 32'd7036;
			58501: outdata = 32'd7035;
			58502: outdata = 32'd7034;
			58503: outdata = 32'd7033;
			58504: outdata = 32'd7032;
			58505: outdata = 32'd7031;
			58506: outdata = 32'd7030;
			58507: outdata = 32'd7029;
			58508: outdata = 32'd7028;
			58509: outdata = 32'd7027;
			58510: outdata = 32'd7026;
			58511: outdata = 32'd7025;
			58512: outdata = 32'd7024;
			58513: outdata = 32'd7023;
			58514: outdata = 32'd7022;
			58515: outdata = 32'd7021;
			58516: outdata = 32'd7020;
			58517: outdata = 32'd7019;
			58518: outdata = 32'd7018;
			58519: outdata = 32'd7017;
			58520: outdata = 32'd7016;
			58521: outdata = 32'd7015;
			58522: outdata = 32'd7014;
			58523: outdata = 32'd7013;
			58524: outdata = 32'd7012;
			58525: outdata = 32'd7011;
			58526: outdata = 32'd7010;
			58527: outdata = 32'd7009;
			58528: outdata = 32'd7008;
			58529: outdata = 32'd7007;
			58530: outdata = 32'd7006;
			58531: outdata = 32'd7005;
			58532: outdata = 32'd7004;
			58533: outdata = 32'd7003;
			58534: outdata = 32'd7002;
			58535: outdata = 32'd7001;
			58536: outdata = 32'd7000;
			58537: outdata = 32'd6999;
			58538: outdata = 32'd6998;
			58539: outdata = 32'd6997;
			58540: outdata = 32'd6996;
			58541: outdata = 32'd6995;
			58542: outdata = 32'd6994;
			58543: outdata = 32'd6993;
			58544: outdata = 32'd6992;
			58545: outdata = 32'd6991;
			58546: outdata = 32'd6990;
			58547: outdata = 32'd6989;
			58548: outdata = 32'd6988;
			58549: outdata = 32'd6987;
			58550: outdata = 32'd6986;
			58551: outdata = 32'd6985;
			58552: outdata = 32'd6984;
			58553: outdata = 32'd6983;
			58554: outdata = 32'd6982;
			58555: outdata = 32'd6981;
			58556: outdata = 32'd6980;
			58557: outdata = 32'd6979;
			58558: outdata = 32'd6978;
			58559: outdata = 32'd6977;
			58560: outdata = 32'd6976;
			58561: outdata = 32'd6975;
			58562: outdata = 32'd6974;
			58563: outdata = 32'd6973;
			58564: outdata = 32'd6972;
			58565: outdata = 32'd6971;
			58566: outdata = 32'd6970;
			58567: outdata = 32'd6969;
			58568: outdata = 32'd6968;
			58569: outdata = 32'd6967;
			58570: outdata = 32'd6966;
			58571: outdata = 32'd6965;
			58572: outdata = 32'd6964;
			58573: outdata = 32'd6963;
			58574: outdata = 32'd6962;
			58575: outdata = 32'd6961;
			58576: outdata = 32'd6960;
			58577: outdata = 32'd6959;
			58578: outdata = 32'd6958;
			58579: outdata = 32'd6957;
			58580: outdata = 32'd6956;
			58581: outdata = 32'd6955;
			58582: outdata = 32'd6954;
			58583: outdata = 32'd6953;
			58584: outdata = 32'd6952;
			58585: outdata = 32'd6951;
			58586: outdata = 32'd6950;
			58587: outdata = 32'd6949;
			58588: outdata = 32'd6948;
			58589: outdata = 32'd6947;
			58590: outdata = 32'd6946;
			58591: outdata = 32'd6945;
			58592: outdata = 32'd6944;
			58593: outdata = 32'd6943;
			58594: outdata = 32'd6942;
			58595: outdata = 32'd6941;
			58596: outdata = 32'd6940;
			58597: outdata = 32'd6939;
			58598: outdata = 32'd6938;
			58599: outdata = 32'd6937;
			58600: outdata = 32'd6936;
			58601: outdata = 32'd6935;
			58602: outdata = 32'd6934;
			58603: outdata = 32'd6933;
			58604: outdata = 32'd6932;
			58605: outdata = 32'd6931;
			58606: outdata = 32'd6930;
			58607: outdata = 32'd6929;
			58608: outdata = 32'd6928;
			58609: outdata = 32'd6927;
			58610: outdata = 32'd6926;
			58611: outdata = 32'd6925;
			58612: outdata = 32'd6924;
			58613: outdata = 32'd6923;
			58614: outdata = 32'd6922;
			58615: outdata = 32'd6921;
			58616: outdata = 32'd6920;
			58617: outdata = 32'd6919;
			58618: outdata = 32'd6918;
			58619: outdata = 32'd6917;
			58620: outdata = 32'd6916;
			58621: outdata = 32'd6915;
			58622: outdata = 32'd6914;
			58623: outdata = 32'd6913;
			58624: outdata = 32'd6912;
			58625: outdata = 32'd6911;
			58626: outdata = 32'd6910;
			58627: outdata = 32'd6909;
			58628: outdata = 32'd6908;
			58629: outdata = 32'd6907;
			58630: outdata = 32'd6906;
			58631: outdata = 32'd6905;
			58632: outdata = 32'd6904;
			58633: outdata = 32'd6903;
			58634: outdata = 32'd6902;
			58635: outdata = 32'd6901;
			58636: outdata = 32'd6900;
			58637: outdata = 32'd6899;
			58638: outdata = 32'd6898;
			58639: outdata = 32'd6897;
			58640: outdata = 32'd6896;
			58641: outdata = 32'd6895;
			58642: outdata = 32'd6894;
			58643: outdata = 32'd6893;
			58644: outdata = 32'd6892;
			58645: outdata = 32'd6891;
			58646: outdata = 32'd6890;
			58647: outdata = 32'd6889;
			58648: outdata = 32'd6888;
			58649: outdata = 32'd6887;
			58650: outdata = 32'd6886;
			58651: outdata = 32'd6885;
			58652: outdata = 32'd6884;
			58653: outdata = 32'd6883;
			58654: outdata = 32'd6882;
			58655: outdata = 32'd6881;
			58656: outdata = 32'd6880;
			58657: outdata = 32'd6879;
			58658: outdata = 32'd6878;
			58659: outdata = 32'd6877;
			58660: outdata = 32'd6876;
			58661: outdata = 32'd6875;
			58662: outdata = 32'd6874;
			58663: outdata = 32'd6873;
			58664: outdata = 32'd6872;
			58665: outdata = 32'd6871;
			58666: outdata = 32'd6870;
			58667: outdata = 32'd6869;
			58668: outdata = 32'd6868;
			58669: outdata = 32'd6867;
			58670: outdata = 32'd6866;
			58671: outdata = 32'd6865;
			58672: outdata = 32'd6864;
			58673: outdata = 32'd6863;
			58674: outdata = 32'd6862;
			58675: outdata = 32'd6861;
			58676: outdata = 32'd6860;
			58677: outdata = 32'd6859;
			58678: outdata = 32'd6858;
			58679: outdata = 32'd6857;
			58680: outdata = 32'd6856;
			58681: outdata = 32'd6855;
			58682: outdata = 32'd6854;
			58683: outdata = 32'd6853;
			58684: outdata = 32'd6852;
			58685: outdata = 32'd6851;
			58686: outdata = 32'd6850;
			58687: outdata = 32'd6849;
			58688: outdata = 32'd6848;
			58689: outdata = 32'd6847;
			58690: outdata = 32'd6846;
			58691: outdata = 32'd6845;
			58692: outdata = 32'd6844;
			58693: outdata = 32'd6843;
			58694: outdata = 32'd6842;
			58695: outdata = 32'd6841;
			58696: outdata = 32'd6840;
			58697: outdata = 32'd6839;
			58698: outdata = 32'd6838;
			58699: outdata = 32'd6837;
			58700: outdata = 32'd6836;
			58701: outdata = 32'd6835;
			58702: outdata = 32'd6834;
			58703: outdata = 32'd6833;
			58704: outdata = 32'd6832;
			58705: outdata = 32'd6831;
			58706: outdata = 32'd6830;
			58707: outdata = 32'd6829;
			58708: outdata = 32'd6828;
			58709: outdata = 32'd6827;
			58710: outdata = 32'd6826;
			58711: outdata = 32'd6825;
			58712: outdata = 32'd6824;
			58713: outdata = 32'd6823;
			58714: outdata = 32'd6822;
			58715: outdata = 32'd6821;
			58716: outdata = 32'd6820;
			58717: outdata = 32'd6819;
			58718: outdata = 32'd6818;
			58719: outdata = 32'd6817;
			58720: outdata = 32'd6816;
			58721: outdata = 32'd6815;
			58722: outdata = 32'd6814;
			58723: outdata = 32'd6813;
			58724: outdata = 32'd6812;
			58725: outdata = 32'd6811;
			58726: outdata = 32'd6810;
			58727: outdata = 32'd6809;
			58728: outdata = 32'd6808;
			58729: outdata = 32'd6807;
			58730: outdata = 32'd6806;
			58731: outdata = 32'd6805;
			58732: outdata = 32'd6804;
			58733: outdata = 32'd6803;
			58734: outdata = 32'd6802;
			58735: outdata = 32'd6801;
			58736: outdata = 32'd6800;
			58737: outdata = 32'd6799;
			58738: outdata = 32'd6798;
			58739: outdata = 32'd6797;
			58740: outdata = 32'd6796;
			58741: outdata = 32'd6795;
			58742: outdata = 32'd6794;
			58743: outdata = 32'd6793;
			58744: outdata = 32'd6792;
			58745: outdata = 32'd6791;
			58746: outdata = 32'd6790;
			58747: outdata = 32'd6789;
			58748: outdata = 32'd6788;
			58749: outdata = 32'd6787;
			58750: outdata = 32'd6786;
			58751: outdata = 32'd6785;
			58752: outdata = 32'd6784;
			58753: outdata = 32'd6783;
			58754: outdata = 32'd6782;
			58755: outdata = 32'd6781;
			58756: outdata = 32'd6780;
			58757: outdata = 32'd6779;
			58758: outdata = 32'd6778;
			58759: outdata = 32'd6777;
			58760: outdata = 32'd6776;
			58761: outdata = 32'd6775;
			58762: outdata = 32'd6774;
			58763: outdata = 32'd6773;
			58764: outdata = 32'd6772;
			58765: outdata = 32'd6771;
			58766: outdata = 32'd6770;
			58767: outdata = 32'd6769;
			58768: outdata = 32'd6768;
			58769: outdata = 32'd6767;
			58770: outdata = 32'd6766;
			58771: outdata = 32'd6765;
			58772: outdata = 32'd6764;
			58773: outdata = 32'd6763;
			58774: outdata = 32'd6762;
			58775: outdata = 32'd6761;
			58776: outdata = 32'd6760;
			58777: outdata = 32'd6759;
			58778: outdata = 32'd6758;
			58779: outdata = 32'd6757;
			58780: outdata = 32'd6756;
			58781: outdata = 32'd6755;
			58782: outdata = 32'd6754;
			58783: outdata = 32'd6753;
			58784: outdata = 32'd6752;
			58785: outdata = 32'd6751;
			58786: outdata = 32'd6750;
			58787: outdata = 32'd6749;
			58788: outdata = 32'd6748;
			58789: outdata = 32'd6747;
			58790: outdata = 32'd6746;
			58791: outdata = 32'd6745;
			58792: outdata = 32'd6744;
			58793: outdata = 32'd6743;
			58794: outdata = 32'd6742;
			58795: outdata = 32'd6741;
			58796: outdata = 32'd6740;
			58797: outdata = 32'd6739;
			58798: outdata = 32'd6738;
			58799: outdata = 32'd6737;
			58800: outdata = 32'd6736;
			58801: outdata = 32'd6735;
			58802: outdata = 32'd6734;
			58803: outdata = 32'd6733;
			58804: outdata = 32'd6732;
			58805: outdata = 32'd6731;
			58806: outdata = 32'd6730;
			58807: outdata = 32'd6729;
			58808: outdata = 32'd6728;
			58809: outdata = 32'd6727;
			58810: outdata = 32'd6726;
			58811: outdata = 32'd6725;
			58812: outdata = 32'd6724;
			58813: outdata = 32'd6723;
			58814: outdata = 32'd6722;
			58815: outdata = 32'd6721;
			58816: outdata = 32'd6720;
			58817: outdata = 32'd6719;
			58818: outdata = 32'd6718;
			58819: outdata = 32'd6717;
			58820: outdata = 32'd6716;
			58821: outdata = 32'd6715;
			58822: outdata = 32'd6714;
			58823: outdata = 32'd6713;
			58824: outdata = 32'd6712;
			58825: outdata = 32'd6711;
			58826: outdata = 32'd6710;
			58827: outdata = 32'd6709;
			58828: outdata = 32'd6708;
			58829: outdata = 32'd6707;
			58830: outdata = 32'd6706;
			58831: outdata = 32'd6705;
			58832: outdata = 32'd6704;
			58833: outdata = 32'd6703;
			58834: outdata = 32'd6702;
			58835: outdata = 32'd6701;
			58836: outdata = 32'd6700;
			58837: outdata = 32'd6699;
			58838: outdata = 32'd6698;
			58839: outdata = 32'd6697;
			58840: outdata = 32'd6696;
			58841: outdata = 32'd6695;
			58842: outdata = 32'd6694;
			58843: outdata = 32'd6693;
			58844: outdata = 32'd6692;
			58845: outdata = 32'd6691;
			58846: outdata = 32'd6690;
			58847: outdata = 32'd6689;
			58848: outdata = 32'd6688;
			58849: outdata = 32'd6687;
			58850: outdata = 32'd6686;
			58851: outdata = 32'd6685;
			58852: outdata = 32'd6684;
			58853: outdata = 32'd6683;
			58854: outdata = 32'd6682;
			58855: outdata = 32'd6681;
			58856: outdata = 32'd6680;
			58857: outdata = 32'd6679;
			58858: outdata = 32'd6678;
			58859: outdata = 32'd6677;
			58860: outdata = 32'd6676;
			58861: outdata = 32'd6675;
			58862: outdata = 32'd6674;
			58863: outdata = 32'd6673;
			58864: outdata = 32'd6672;
			58865: outdata = 32'd6671;
			58866: outdata = 32'd6670;
			58867: outdata = 32'd6669;
			58868: outdata = 32'd6668;
			58869: outdata = 32'd6667;
			58870: outdata = 32'd6666;
			58871: outdata = 32'd6665;
			58872: outdata = 32'd6664;
			58873: outdata = 32'd6663;
			58874: outdata = 32'd6662;
			58875: outdata = 32'd6661;
			58876: outdata = 32'd6660;
			58877: outdata = 32'd6659;
			58878: outdata = 32'd6658;
			58879: outdata = 32'd6657;
			58880: outdata = 32'd6656;
			58881: outdata = 32'd6655;
			58882: outdata = 32'd6654;
			58883: outdata = 32'd6653;
			58884: outdata = 32'd6652;
			58885: outdata = 32'd6651;
			58886: outdata = 32'd6650;
			58887: outdata = 32'd6649;
			58888: outdata = 32'd6648;
			58889: outdata = 32'd6647;
			58890: outdata = 32'd6646;
			58891: outdata = 32'd6645;
			58892: outdata = 32'd6644;
			58893: outdata = 32'd6643;
			58894: outdata = 32'd6642;
			58895: outdata = 32'd6641;
			58896: outdata = 32'd6640;
			58897: outdata = 32'd6639;
			58898: outdata = 32'd6638;
			58899: outdata = 32'd6637;
			58900: outdata = 32'd6636;
			58901: outdata = 32'd6635;
			58902: outdata = 32'd6634;
			58903: outdata = 32'd6633;
			58904: outdata = 32'd6632;
			58905: outdata = 32'd6631;
			58906: outdata = 32'd6630;
			58907: outdata = 32'd6629;
			58908: outdata = 32'd6628;
			58909: outdata = 32'd6627;
			58910: outdata = 32'd6626;
			58911: outdata = 32'd6625;
			58912: outdata = 32'd6624;
			58913: outdata = 32'd6623;
			58914: outdata = 32'd6622;
			58915: outdata = 32'd6621;
			58916: outdata = 32'd6620;
			58917: outdata = 32'd6619;
			58918: outdata = 32'd6618;
			58919: outdata = 32'd6617;
			58920: outdata = 32'd6616;
			58921: outdata = 32'd6615;
			58922: outdata = 32'd6614;
			58923: outdata = 32'd6613;
			58924: outdata = 32'd6612;
			58925: outdata = 32'd6611;
			58926: outdata = 32'd6610;
			58927: outdata = 32'd6609;
			58928: outdata = 32'd6608;
			58929: outdata = 32'd6607;
			58930: outdata = 32'd6606;
			58931: outdata = 32'd6605;
			58932: outdata = 32'd6604;
			58933: outdata = 32'd6603;
			58934: outdata = 32'd6602;
			58935: outdata = 32'd6601;
			58936: outdata = 32'd6600;
			58937: outdata = 32'd6599;
			58938: outdata = 32'd6598;
			58939: outdata = 32'd6597;
			58940: outdata = 32'd6596;
			58941: outdata = 32'd6595;
			58942: outdata = 32'd6594;
			58943: outdata = 32'd6593;
			58944: outdata = 32'd6592;
			58945: outdata = 32'd6591;
			58946: outdata = 32'd6590;
			58947: outdata = 32'd6589;
			58948: outdata = 32'd6588;
			58949: outdata = 32'd6587;
			58950: outdata = 32'd6586;
			58951: outdata = 32'd6585;
			58952: outdata = 32'd6584;
			58953: outdata = 32'd6583;
			58954: outdata = 32'd6582;
			58955: outdata = 32'd6581;
			58956: outdata = 32'd6580;
			58957: outdata = 32'd6579;
			58958: outdata = 32'd6578;
			58959: outdata = 32'd6577;
			58960: outdata = 32'd6576;
			58961: outdata = 32'd6575;
			58962: outdata = 32'd6574;
			58963: outdata = 32'd6573;
			58964: outdata = 32'd6572;
			58965: outdata = 32'd6571;
			58966: outdata = 32'd6570;
			58967: outdata = 32'd6569;
			58968: outdata = 32'd6568;
			58969: outdata = 32'd6567;
			58970: outdata = 32'd6566;
			58971: outdata = 32'd6565;
			58972: outdata = 32'd6564;
			58973: outdata = 32'd6563;
			58974: outdata = 32'd6562;
			58975: outdata = 32'd6561;
			58976: outdata = 32'd6560;
			58977: outdata = 32'd6559;
			58978: outdata = 32'd6558;
			58979: outdata = 32'd6557;
			58980: outdata = 32'd6556;
			58981: outdata = 32'd6555;
			58982: outdata = 32'd6554;
			58983: outdata = 32'd6553;
			58984: outdata = 32'd6552;
			58985: outdata = 32'd6551;
			58986: outdata = 32'd6550;
			58987: outdata = 32'd6549;
			58988: outdata = 32'd6548;
			58989: outdata = 32'd6547;
			58990: outdata = 32'd6546;
			58991: outdata = 32'd6545;
			58992: outdata = 32'd6544;
			58993: outdata = 32'd6543;
			58994: outdata = 32'd6542;
			58995: outdata = 32'd6541;
			58996: outdata = 32'd6540;
			58997: outdata = 32'd6539;
			58998: outdata = 32'd6538;
			58999: outdata = 32'd6537;
			59000: outdata = 32'd6536;
			59001: outdata = 32'd6535;
			59002: outdata = 32'd6534;
			59003: outdata = 32'd6533;
			59004: outdata = 32'd6532;
			59005: outdata = 32'd6531;
			59006: outdata = 32'd6530;
			59007: outdata = 32'd6529;
			59008: outdata = 32'd6528;
			59009: outdata = 32'd6527;
			59010: outdata = 32'd6526;
			59011: outdata = 32'd6525;
			59012: outdata = 32'd6524;
			59013: outdata = 32'd6523;
			59014: outdata = 32'd6522;
			59015: outdata = 32'd6521;
			59016: outdata = 32'd6520;
			59017: outdata = 32'd6519;
			59018: outdata = 32'd6518;
			59019: outdata = 32'd6517;
			59020: outdata = 32'd6516;
			59021: outdata = 32'd6515;
			59022: outdata = 32'd6514;
			59023: outdata = 32'd6513;
			59024: outdata = 32'd6512;
			59025: outdata = 32'd6511;
			59026: outdata = 32'd6510;
			59027: outdata = 32'd6509;
			59028: outdata = 32'd6508;
			59029: outdata = 32'd6507;
			59030: outdata = 32'd6506;
			59031: outdata = 32'd6505;
			59032: outdata = 32'd6504;
			59033: outdata = 32'd6503;
			59034: outdata = 32'd6502;
			59035: outdata = 32'd6501;
			59036: outdata = 32'd6500;
			59037: outdata = 32'd6499;
			59038: outdata = 32'd6498;
			59039: outdata = 32'd6497;
			59040: outdata = 32'd6496;
			59041: outdata = 32'd6495;
			59042: outdata = 32'd6494;
			59043: outdata = 32'd6493;
			59044: outdata = 32'd6492;
			59045: outdata = 32'd6491;
			59046: outdata = 32'd6490;
			59047: outdata = 32'd6489;
			59048: outdata = 32'd6488;
			59049: outdata = 32'd6487;
			59050: outdata = 32'd6486;
			59051: outdata = 32'd6485;
			59052: outdata = 32'd6484;
			59053: outdata = 32'd6483;
			59054: outdata = 32'd6482;
			59055: outdata = 32'd6481;
			59056: outdata = 32'd6480;
			59057: outdata = 32'd6479;
			59058: outdata = 32'd6478;
			59059: outdata = 32'd6477;
			59060: outdata = 32'd6476;
			59061: outdata = 32'd6475;
			59062: outdata = 32'd6474;
			59063: outdata = 32'd6473;
			59064: outdata = 32'd6472;
			59065: outdata = 32'd6471;
			59066: outdata = 32'd6470;
			59067: outdata = 32'd6469;
			59068: outdata = 32'd6468;
			59069: outdata = 32'd6467;
			59070: outdata = 32'd6466;
			59071: outdata = 32'd6465;
			59072: outdata = 32'd6464;
			59073: outdata = 32'd6463;
			59074: outdata = 32'd6462;
			59075: outdata = 32'd6461;
			59076: outdata = 32'd6460;
			59077: outdata = 32'd6459;
			59078: outdata = 32'd6458;
			59079: outdata = 32'd6457;
			59080: outdata = 32'd6456;
			59081: outdata = 32'd6455;
			59082: outdata = 32'd6454;
			59083: outdata = 32'd6453;
			59084: outdata = 32'd6452;
			59085: outdata = 32'd6451;
			59086: outdata = 32'd6450;
			59087: outdata = 32'd6449;
			59088: outdata = 32'd6448;
			59089: outdata = 32'd6447;
			59090: outdata = 32'd6446;
			59091: outdata = 32'd6445;
			59092: outdata = 32'd6444;
			59093: outdata = 32'd6443;
			59094: outdata = 32'd6442;
			59095: outdata = 32'd6441;
			59096: outdata = 32'd6440;
			59097: outdata = 32'd6439;
			59098: outdata = 32'd6438;
			59099: outdata = 32'd6437;
			59100: outdata = 32'd6436;
			59101: outdata = 32'd6435;
			59102: outdata = 32'd6434;
			59103: outdata = 32'd6433;
			59104: outdata = 32'd6432;
			59105: outdata = 32'd6431;
			59106: outdata = 32'd6430;
			59107: outdata = 32'd6429;
			59108: outdata = 32'd6428;
			59109: outdata = 32'd6427;
			59110: outdata = 32'd6426;
			59111: outdata = 32'd6425;
			59112: outdata = 32'd6424;
			59113: outdata = 32'd6423;
			59114: outdata = 32'd6422;
			59115: outdata = 32'd6421;
			59116: outdata = 32'd6420;
			59117: outdata = 32'd6419;
			59118: outdata = 32'd6418;
			59119: outdata = 32'd6417;
			59120: outdata = 32'd6416;
			59121: outdata = 32'd6415;
			59122: outdata = 32'd6414;
			59123: outdata = 32'd6413;
			59124: outdata = 32'd6412;
			59125: outdata = 32'd6411;
			59126: outdata = 32'd6410;
			59127: outdata = 32'd6409;
			59128: outdata = 32'd6408;
			59129: outdata = 32'd6407;
			59130: outdata = 32'd6406;
			59131: outdata = 32'd6405;
			59132: outdata = 32'd6404;
			59133: outdata = 32'd6403;
			59134: outdata = 32'd6402;
			59135: outdata = 32'd6401;
			59136: outdata = 32'd6400;
			59137: outdata = 32'd6399;
			59138: outdata = 32'd6398;
			59139: outdata = 32'd6397;
			59140: outdata = 32'd6396;
			59141: outdata = 32'd6395;
			59142: outdata = 32'd6394;
			59143: outdata = 32'd6393;
			59144: outdata = 32'd6392;
			59145: outdata = 32'd6391;
			59146: outdata = 32'd6390;
			59147: outdata = 32'd6389;
			59148: outdata = 32'd6388;
			59149: outdata = 32'd6387;
			59150: outdata = 32'd6386;
			59151: outdata = 32'd6385;
			59152: outdata = 32'd6384;
			59153: outdata = 32'd6383;
			59154: outdata = 32'd6382;
			59155: outdata = 32'd6381;
			59156: outdata = 32'd6380;
			59157: outdata = 32'd6379;
			59158: outdata = 32'd6378;
			59159: outdata = 32'd6377;
			59160: outdata = 32'd6376;
			59161: outdata = 32'd6375;
			59162: outdata = 32'd6374;
			59163: outdata = 32'd6373;
			59164: outdata = 32'd6372;
			59165: outdata = 32'd6371;
			59166: outdata = 32'd6370;
			59167: outdata = 32'd6369;
			59168: outdata = 32'd6368;
			59169: outdata = 32'd6367;
			59170: outdata = 32'd6366;
			59171: outdata = 32'd6365;
			59172: outdata = 32'd6364;
			59173: outdata = 32'd6363;
			59174: outdata = 32'd6362;
			59175: outdata = 32'd6361;
			59176: outdata = 32'd6360;
			59177: outdata = 32'd6359;
			59178: outdata = 32'd6358;
			59179: outdata = 32'd6357;
			59180: outdata = 32'd6356;
			59181: outdata = 32'd6355;
			59182: outdata = 32'd6354;
			59183: outdata = 32'd6353;
			59184: outdata = 32'd6352;
			59185: outdata = 32'd6351;
			59186: outdata = 32'd6350;
			59187: outdata = 32'd6349;
			59188: outdata = 32'd6348;
			59189: outdata = 32'd6347;
			59190: outdata = 32'd6346;
			59191: outdata = 32'd6345;
			59192: outdata = 32'd6344;
			59193: outdata = 32'd6343;
			59194: outdata = 32'd6342;
			59195: outdata = 32'd6341;
			59196: outdata = 32'd6340;
			59197: outdata = 32'd6339;
			59198: outdata = 32'd6338;
			59199: outdata = 32'd6337;
			59200: outdata = 32'd6336;
			59201: outdata = 32'd6335;
			59202: outdata = 32'd6334;
			59203: outdata = 32'd6333;
			59204: outdata = 32'd6332;
			59205: outdata = 32'd6331;
			59206: outdata = 32'd6330;
			59207: outdata = 32'd6329;
			59208: outdata = 32'd6328;
			59209: outdata = 32'd6327;
			59210: outdata = 32'd6326;
			59211: outdata = 32'd6325;
			59212: outdata = 32'd6324;
			59213: outdata = 32'd6323;
			59214: outdata = 32'd6322;
			59215: outdata = 32'd6321;
			59216: outdata = 32'd6320;
			59217: outdata = 32'd6319;
			59218: outdata = 32'd6318;
			59219: outdata = 32'd6317;
			59220: outdata = 32'd6316;
			59221: outdata = 32'd6315;
			59222: outdata = 32'd6314;
			59223: outdata = 32'd6313;
			59224: outdata = 32'd6312;
			59225: outdata = 32'd6311;
			59226: outdata = 32'd6310;
			59227: outdata = 32'd6309;
			59228: outdata = 32'd6308;
			59229: outdata = 32'd6307;
			59230: outdata = 32'd6306;
			59231: outdata = 32'd6305;
			59232: outdata = 32'd6304;
			59233: outdata = 32'd6303;
			59234: outdata = 32'd6302;
			59235: outdata = 32'd6301;
			59236: outdata = 32'd6300;
			59237: outdata = 32'd6299;
			59238: outdata = 32'd6298;
			59239: outdata = 32'd6297;
			59240: outdata = 32'd6296;
			59241: outdata = 32'd6295;
			59242: outdata = 32'd6294;
			59243: outdata = 32'd6293;
			59244: outdata = 32'd6292;
			59245: outdata = 32'd6291;
			59246: outdata = 32'd6290;
			59247: outdata = 32'd6289;
			59248: outdata = 32'd6288;
			59249: outdata = 32'd6287;
			59250: outdata = 32'd6286;
			59251: outdata = 32'd6285;
			59252: outdata = 32'd6284;
			59253: outdata = 32'd6283;
			59254: outdata = 32'd6282;
			59255: outdata = 32'd6281;
			59256: outdata = 32'd6280;
			59257: outdata = 32'd6279;
			59258: outdata = 32'd6278;
			59259: outdata = 32'd6277;
			59260: outdata = 32'd6276;
			59261: outdata = 32'd6275;
			59262: outdata = 32'd6274;
			59263: outdata = 32'd6273;
			59264: outdata = 32'd6272;
			59265: outdata = 32'd6271;
			59266: outdata = 32'd6270;
			59267: outdata = 32'd6269;
			59268: outdata = 32'd6268;
			59269: outdata = 32'd6267;
			59270: outdata = 32'd6266;
			59271: outdata = 32'd6265;
			59272: outdata = 32'd6264;
			59273: outdata = 32'd6263;
			59274: outdata = 32'd6262;
			59275: outdata = 32'd6261;
			59276: outdata = 32'd6260;
			59277: outdata = 32'd6259;
			59278: outdata = 32'd6258;
			59279: outdata = 32'd6257;
			59280: outdata = 32'd6256;
			59281: outdata = 32'd6255;
			59282: outdata = 32'd6254;
			59283: outdata = 32'd6253;
			59284: outdata = 32'd6252;
			59285: outdata = 32'd6251;
			59286: outdata = 32'd6250;
			59287: outdata = 32'd6249;
			59288: outdata = 32'd6248;
			59289: outdata = 32'd6247;
			59290: outdata = 32'd6246;
			59291: outdata = 32'd6245;
			59292: outdata = 32'd6244;
			59293: outdata = 32'd6243;
			59294: outdata = 32'd6242;
			59295: outdata = 32'd6241;
			59296: outdata = 32'd6240;
			59297: outdata = 32'd6239;
			59298: outdata = 32'd6238;
			59299: outdata = 32'd6237;
			59300: outdata = 32'd6236;
			59301: outdata = 32'd6235;
			59302: outdata = 32'd6234;
			59303: outdata = 32'd6233;
			59304: outdata = 32'd6232;
			59305: outdata = 32'd6231;
			59306: outdata = 32'd6230;
			59307: outdata = 32'd6229;
			59308: outdata = 32'd6228;
			59309: outdata = 32'd6227;
			59310: outdata = 32'd6226;
			59311: outdata = 32'd6225;
			59312: outdata = 32'd6224;
			59313: outdata = 32'd6223;
			59314: outdata = 32'd6222;
			59315: outdata = 32'd6221;
			59316: outdata = 32'd6220;
			59317: outdata = 32'd6219;
			59318: outdata = 32'd6218;
			59319: outdata = 32'd6217;
			59320: outdata = 32'd6216;
			59321: outdata = 32'd6215;
			59322: outdata = 32'd6214;
			59323: outdata = 32'd6213;
			59324: outdata = 32'd6212;
			59325: outdata = 32'd6211;
			59326: outdata = 32'd6210;
			59327: outdata = 32'd6209;
			59328: outdata = 32'd6208;
			59329: outdata = 32'd6207;
			59330: outdata = 32'd6206;
			59331: outdata = 32'd6205;
			59332: outdata = 32'd6204;
			59333: outdata = 32'd6203;
			59334: outdata = 32'd6202;
			59335: outdata = 32'd6201;
			59336: outdata = 32'd6200;
			59337: outdata = 32'd6199;
			59338: outdata = 32'd6198;
			59339: outdata = 32'd6197;
			59340: outdata = 32'd6196;
			59341: outdata = 32'd6195;
			59342: outdata = 32'd6194;
			59343: outdata = 32'd6193;
			59344: outdata = 32'd6192;
			59345: outdata = 32'd6191;
			59346: outdata = 32'd6190;
			59347: outdata = 32'd6189;
			59348: outdata = 32'd6188;
			59349: outdata = 32'd6187;
			59350: outdata = 32'd6186;
			59351: outdata = 32'd6185;
			59352: outdata = 32'd6184;
			59353: outdata = 32'd6183;
			59354: outdata = 32'd6182;
			59355: outdata = 32'd6181;
			59356: outdata = 32'd6180;
			59357: outdata = 32'd6179;
			59358: outdata = 32'd6178;
			59359: outdata = 32'd6177;
			59360: outdata = 32'd6176;
			59361: outdata = 32'd6175;
			59362: outdata = 32'd6174;
			59363: outdata = 32'd6173;
			59364: outdata = 32'd6172;
			59365: outdata = 32'd6171;
			59366: outdata = 32'd6170;
			59367: outdata = 32'd6169;
			59368: outdata = 32'd6168;
			59369: outdata = 32'd6167;
			59370: outdata = 32'd6166;
			59371: outdata = 32'd6165;
			59372: outdata = 32'd6164;
			59373: outdata = 32'd6163;
			59374: outdata = 32'd6162;
			59375: outdata = 32'd6161;
			59376: outdata = 32'd6160;
			59377: outdata = 32'd6159;
			59378: outdata = 32'd6158;
			59379: outdata = 32'd6157;
			59380: outdata = 32'd6156;
			59381: outdata = 32'd6155;
			59382: outdata = 32'd6154;
			59383: outdata = 32'd6153;
			59384: outdata = 32'd6152;
			59385: outdata = 32'd6151;
			59386: outdata = 32'd6150;
			59387: outdata = 32'd6149;
			59388: outdata = 32'd6148;
			59389: outdata = 32'd6147;
			59390: outdata = 32'd6146;
			59391: outdata = 32'd6145;
			59392: outdata = 32'd6144;
			59393: outdata = 32'd6143;
			59394: outdata = 32'd6142;
			59395: outdata = 32'd6141;
			59396: outdata = 32'd6140;
			59397: outdata = 32'd6139;
			59398: outdata = 32'd6138;
			59399: outdata = 32'd6137;
			59400: outdata = 32'd6136;
			59401: outdata = 32'd6135;
			59402: outdata = 32'd6134;
			59403: outdata = 32'd6133;
			59404: outdata = 32'd6132;
			59405: outdata = 32'd6131;
			59406: outdata = 32'd6130;
			59407: outdata = 32'd6129;
			59408: outdata = 32'd6128;
			59409: outdata = 32'd6127;
			59410: outdata = 32'd6126;
			59411: outdata = 32'd6125;
			59412: outdata = 32'd6124;
			59413: outdata = 32'd6123;
			59414: outdata = 32'd6122;
			59415: outdata = 32'd6121;
			59416: outdata = 32'd6120;
			59417: outdata = 32'd6119;
			59418: outdata = 32'd6118;
			59419: outdata = 32'd6117;
			59420: outdata = 32'd6116;
			59421: outdata = 32'd6115;
			59422: outdata = 32'd6114;
			59423: outdata = 32'd6113;
			59424: outdata = 32'd6112;
			59425: outdata = 32'd6111;
			59426: outdata = 32'd6110;
			59427: outdata = 32'd6109;
			59428: outdata = 32'd6108;
			59429: outdata = 32'd6107;
			59430: outdata = 32'd6106;
			59431: outdata = 32'd6105;
			59432: outdata = 32'd6104;
			59433: outdata = 32'd6103;
			59434: outdata = 32'd6102;
			59435: outdata = 32'd6101;
			59436: outdata = 32'd6100;
			59437: outdata = 32'd6099;
			59438: outdata = 32'd6098;
			59439: outdata = 32'd6097;
			59440: outdata = 32'd6096;
			59441: outdata = 32'd6095;
			59442: outdata = 32'd6094;
			59443: outdata = 32'd6093;
			59444: outdata = 32'd6092;
			59445: outdata = 32'd6091;
			59446: outdata = 32'd6090;
			59447: outdata = 32'd6089;
			59448: outdata = 32'd6088;
			59449: outdata = 32'd6087;
			59450: outdata = 32'd6086;
			59451: outdata = 32'd6085;
			59452: outdata = 32'd6084;
			59453: outdata = 32'd6083;
			59454: outdata = 32'd6082;
			59455: outdata = 32'd6081;
			59456: outdata = 32'd6080;
			59457: outdata = 32'd6079;
			59458: outdata = 32'd6078;
			59459: outdata = 32'd6077;
			59460: outdata = 32'd6076;
			59461: outdata = 32'd6075;
			59462: outdata = 32'd6074;
			59463: outdata = 32'd6073;
			59464: outdata = 32'd6072;
			59465: outdata = 32'd6071;
			59466: outdata = 32'd6070;
			59467: outdata = 32'd6069;
			59468: outdata = 32'd6068;
			59469: outdata = 32'd6067;
			59470: outdata = 32'd6066;
			59471: outdata = 32'd6065;
			59472: outdata = 32'd6064;
			59473: outdata = 32'd6063;
			59474: outdata = 32'd6062;
			59475: outdata = 32'd6061;
			59476: outdata = 32'd6060;
			59477: outdata = 32'd6059;
			59478: outdata = 32'd6058;
			59479: outdata = 32'd6057;
			59480: outdata = 32'd6056;
			59481: outdata = 32'd6055;
			59482: outdata = 32'd6054;
			59483: outdata = 32'd6053;
			59484: outdata = 32'd6052;
			59485: outdata = 32'd6051;
			59486: outdata = 32'd6050;
			59487: outdata = 32'd6049;
			59488: outdata = 32'd6048;
			59489: outdata = 32'd6047;
			59490: outdata = 32'd6046;
			59491: outdata = 32'd6045;
			59492: outdata = 32'd6044;
			59493: outdata = 32'd6043;
			59494: outdata = 32'd6042;
			59495: outdata = 32'd6041;
			59496: outdata = 32'd6040;
			59497: outdata = 32'd6039;
			59498: outdata = 32'd6038;
			59499: outdata = 32'd6037;
			59500: outdata = 32'd6036;
			59501: outdata = 32'd6035;
			59502: outdata = 32'd6034;
			59503: outdata = 32'd6033;
			59504: outdata = 32'd6032;
			59505: outdata = 32'd6031;
			59506: outdata = 32'd6030;
			59507: outdata = 32'd6029;
			59508: outdata = 32'd6028;
			59509: outdata = 32'd6027;
			59510: outdata = 32'd6026;
			59511: outdata = 32'd6025;
			59512: outdata = 32'd6024;
			59513: outdata = 32'd6023;
			59514: outdata = 32'd6022;
			59515: outdata = 32'd6021;
			59516: outdata = 32'd6020;
			59517: outdata = 32'd6019;
			59518: outdata = 32'd6018;
			59519: outdata = 32'd6017;
			59520: outdata = 32'd6016;
			59521: outdata = 32'd6015;
			59522: outdata = 32'd6014;
			59523: outdata = 32'd6013;
			59524: outdata = 32'd6012;
			59525: outdata = 32'd6011;
			59526: outdata = 32'd6010;
			59527: outdata = 32'd6009;
			59528: outdata = 32'd6008;
			59529: outdata = 32'd6007;
			59530: outdata = 32'd6006;
			59531: outdata = 32'd6005;
			59532: outdata = 32'd6004;
			59533: outdata = 32'd6003;
			59534: outdata = 32'd6002;
			59535: outdata = 32'd6001;
			59536: outdata = 32'd6000;
			59537: outdata = 32'd5999;
			59538: outdata = 32'd5998;
			59539: outdata = 32'd5997;
			59540: outdata = 32'd5996;
			59541: outdata = 32'd5995;
			59542: outdata = 32'd5994;
			59543: outdata = 32'd5993;
			59544: outdata = 32'd5992;
			59545: outdata = 32'd5991;
			59546: outdata = 32'd5990;
			59547: outdata = 32'd5989;
			59548: outdata = 32'd5988;
			59549: outdata = 32'd5987;
			59550: outdata = 32'd5986;
			59551: outdata = 32'd5985;
			59552: outdata = 32'd5984;
			59553: outdata = 32'd5983;
			59554: outdata = 32'd5982;
			59555: outdata = 32'd5981;
			59556: outdata = 32'd5980;
			59557: outdata = 32'd5979;
			59558: outdata = 32'd5978;
			59559: outdata = 32'd5977;
			59560: outdata = 32'd5976;
			59561: outdata = 32'd5975;
			59562: outdata = 32'd5974;
			59563: outdata = 32'd5973;
			59564: outdata = 32'd5972;
			59565: outdata = 32'd5971;
			59566: outdata = 32'd5970;
			59567: outdata = 32'd5969;
			59568: outdata = 32'd5968;
			59569: outdata = 32'd5967;
			59570: outdata = 32'd5966;
			59571: outdata = 32'd5965;
			59572: outdata = 32'd5964;
			59573: outdata = 32'd5963;
			59574: outdata = 32'd5962;
			59575: outdata = 32'd5961;
			59576: outdata = 32'd5960;
			59577: outdata = 32'd5959;
			59578: outdata = 32'd5958;
			59579: outdata = 32'd5957;
			59580: outdata = 32'd5956;
			59581: outdata = 32'd5955;
			59582: outdata = 32'd5954;
			59583: outdata = 32'd5953;
			59584: outdata = 32'd5952;
			59585: outdata = 32'd5951;
			59586: outdata = 32'd5950;
			59587: outdata = 32'd5949;
			59588: outdata = 32'd5948;
			59589: outdata = 32'd5947;
			59590: outdata = 32'd5946;
			59591: outdata = 32'd5945;
			59592: outdata = 32'd5944;
			59593: outdata = 32'd5943;
			59594: outdata = 32'd5942;
			59595: outdata = 32'd5941;
			59596: outdata = 32'd5940;
			59597: outdata = 32'd5939;
			59598: outdata = 32'd5938;
			59599: outdata = 32'd5937;
			59600: outdata = 32'd5936;
			59601: outdata = 32'd5935;
			59602: outdata = 32'd5934;
			59603: outdata = 32'd5933;
			59604: outdata = 32'd5932;
			59605: outdata = 32'd5931;
			59606: outdata = 32'd5930;
			59607: outdata = 32'd5929;
			59608: outdata = 32'd5928;
			59609: outdata = 32'd5927;
			59610: outdata = 32'd5926;
			59611: outdata = 32'd5925;
			59612: outdata = 32'd5924;
			59613: outdata = 32'd5923;
			59614: outdata = 32'd5922;
			59615: outdata = 32'd5921;
			59616: outdata = 32'd5920;
			59617: outdata = 32'd5919;
			59618: outdata = 32'd5918;
			59619: outdata = 32'd5917;
			59620: outdata = 32'd5916;
			59621: outdata = 32'd5915;
			59622: outdata = 32'd5914;
			59623: outdata = 32'd5913;
			59624: outdata = 32'd5912;
			59625: outdata = 32'd5911;
			59626: outdata = 32'd5910;
			59627: outdata = 32'd5909;
			59628: outdata = 32'd5908;
			59629: outdata = 32'd5907;
			59630: outdata = 32'd5906;
			59631: outdata = 32'd5905;
			59632: outdata = 32'd5904;
			59633: outdata = 32'd5903;
			59634: outdata = 32'd5902;
			59635: outdata = 32'd5901;
			59636: outdata = 32'd5900;
			59637: outdata = 32'd5899;
			59638: outdata = 32'd5898;
			59639: outdata = 32'd5897;
			59640: outdata = 32'd5896;
			59641: outdata = 32'd5895;
			59642: outdata = 32'd5894;
			59643: outdata = 32'd5893;
			59644: outdata = 32'd5892;
			59645: outdata = 32'd5891;
			59646: outdata = 32'd5890;
			59647: outdata = 32'd5889;
			59648: outdata = 32'd5888;
			59649: outdata = 32'd5887;
			59650: outdata = 32'd5886;
			59651: outdata = 32'd5885;
			59652: outdata = 32'd5884;
			59653: outdata = 32'd5883;
			59654: outdata = 32'd5882;
			59655: outdata = 32'd5881;
			59656: outdata = 32'd5880;
			59657: outdata = 32'd5879;
			59658: outdata = 32'd5878;
			59659: outdata = 32'd5877;
			59660: outdata = 32'd5876;
			59661: outdata = 32'd5875;
			59662: outdata = 32'd5874;
			59663: outdata = 32'd5873;
			59664: outdata = 32'd5872;
			59665: outdata = 32'd5871;
			59666: outdata = 32'd5870;
			59667: outdata = 32'd5869;
			59668: outdata = 32'd5868;
			59669: outdata = 32'd5867;
			59670: outdata = 32'd5866;
			59671: outdata = 32'd5865;
			59672: outdata = 32'd5864;
			59673: outdata = 32'd5863;
			59674: outdata = 32'd5862;
			59675: outdata = 32'd5861;
			59676: outdata = 32'd5860;
			59677: outdata = 32'd5859;
			59678: outdata = 32'd5858;
			59679: outdata = 32'd5857;
			59680: outdata = 32'd5856;
			59681: outdata = 32'd5855;
			59682: outdata = 32'd5854;
			59683: outdata = 32'd5853;
			59684: outdata = 32'd5852;
			59685: outdata = 32'd5851;
			59686: outdata = 32'd5850;
			59687: outdata = 32'd5849;
			59688: outdata = 32'd5848;
			59689: outdata = 32'd5847;
			59690: outdata = 32'd5846;
			59691: outdata = 32'd5845;
			59692: outdata = 32'd5844;
			59693: outdata = 32'd5843;
			59694: outdata = 32'd5842;
			59695: outdata = 32'd5841;
			59696: outdata = 32'd5840;
			59697: outdata = 32'd5839;
			59698: outdata = 32'd5838;
			59699: outdata = 32'd5837;
			59700: outdata = 32'd5836;
			59701: outdata = 32'd5835;
			59702: outdata = 32'd5834;
			59703: outdata = 32'd5833;
			59704: outdata = 32'd5832;
			59705: outdata = 32'd5831;
			59706: outdata = 32'd5830;
			59707: outdata = 32'd5829;
			59708: outdata = 32'd5828;
			59709: outdata = 32'd5827;
			59710: outdata = 32'd5826;
			59711: outdata = 32'd5825;
			59712: outdata = 32'd5824;
			59713: outdata = 32'd5823;
			59714: outdata = 32'd5822;
			59715: outdata = 32'd5821;
			59716: outdata = 32'd5820;
			59717: outdata = 32'd5819;
			59718: outdata = 32'd5818;
			59719: outdata = 32'd5817;
			59720: outdata = 32'd5816;
			59721: outdata = 32'd5815;
			59722: outdata = 32'd5814;
			59723: outdata = 32'd5813;
			59724: outdata = 32'd5812;
			59725: outdata = 32'd5811;
			59726: outdata = 32'd5810;
			59727: outdata = 32'd5809;
			59728: outdata = 32'd5808;
			59729: outdata = 32'd5807;
			59730: outdata = 32'd5806;
			59731: outdata = 32'd5805;
			59732: outdata = 32'd5804;
			59733: outdata = 32'd5803;
			59734: outdata = 32'd5802;
			59735: outdata = 32'd5801;
			59736: outdata = 32'd5800;
			59737: outdata = 32'd5799;
			59738: outdata = 32'd5798;
			59739: outdata = 32'd5797;
			59740: outdata = 32'd5796;
			59741: outdata = 32'd5795;
			59742: outdata = 32'd5794;
			59743: outdata = 32'd5793;
			59744: outdata = 32'd5792;
			59745: outdata = 32'd5791;
			59746: outdata = 32'd5790;
			59747: outdata = 32'd5789;
			59748: outdata = 32'd5788;
			59749: outdata = 32'd5787;
			59750: outdata = 32'd5786;
			59751: outdata = 32'd5785;
			59752: outdata = 32'd5784;
			59753: outdata = 32'd5783;
			59754: outdata = 32'd5782;
			59755: outdata = 32'd5781;
			59756: outdata = 32'd5780;
			59757: outdata = 32'd5779;
			59758: outdata = 32'd5778;
			59759: outdata = 32'd5777;
			59760: outdata = 32'd5776;
			59761: outdata = 32'd5775;
			59762: outdata = 32'd5774;
			59763: outdata = 32'd5773;
			59764: outdata = 32'd5772;
			59765: outdata = 32'd5771;
			59766: outdata = 32'd5770;
			59767: outdata = 32'd5769;
			59768: outdata = 32'd5768;
			59769: outdata = 32'd5767;
			59770: outdata = 32'd5766;
			59771: outdata = 32'd5765;
			59772: outdata = 32'd5764;
			59773: outdata = 32'd5763;
			59774: outdata = 32'd5762;
			59775: outdata = 32'd5761;
			59776: outdata = 32'd5760;
			59777: outdata = 32'd5759;
			59778: outdata = 32'd5758;
			59779: outdata = 32'd5757;
			59780: outdata = 32'd5756;
			59781: outdata = 32'd5755;
			59782: outdata = 32'd5754;
			59783: outdata = 32'd5753;
			59784: outdata = 32'd5752;
			59785: outdata = 32'd5751;
			59786: outdata = 32'd5750;
			59787: outdata = 32'd5749;
			59788: outdata = 32'd5748;
			59789: outdata = 32'd5747;
			59790: outdata = 32'd5746;
			59791: outdata = 32'd5745;
			59792: outdata = 32'd5744;
			59793: outdata = 32'd5743;
			59794: outdata = 32'd5742;
			59795: outdata = 32'd5741;
			59796: outdata = 32'd5740;
			59797: outdata = 32'd5739;
			59798: outdata = 32'd5738;
			59799: outdata = 32'd5737;
			59800: outdata = 32'd5736;
			59801: outdata = 32'd5735;
			59802: outdata = 32'd5734;
			59803: outdata = 32'd5733;
			59804: outdata = 32'd5732;
			59805: outdata = 32'd5731;
			59806: outdata = 32'd5730;
			59807: outdata = 32'd5729;
			59808: outdata = 32'd5728;
			59809: outdata = 32'd5727;
			59810: outdata = 32'd5726;
			59811: outdata = 32'd5725;
			59812: outdata = 32'd5724;
			59813: outdata = 32'd5723;
			59814: outdata = 32'd5722;
			59815: outdata = 32'd5721;
			59816: outdata = 32'd5720;
			59817: outdata = 32'd5719;
			59818: outdata = 32'd5718;
			59819: outdata = 32'd5717;
			59820: outdata = 32'd5716;
			59821: outdata = 32'd5715;
			59822: outdata = 32'd5714;
			59823: outdata = 32'd5713;
			59824: outdata = 32'd5712;
			59825: outdata = 32'd5711;
			59826: outdata = 32'd5710;
			59827: outdata = 32'd5709;
			59828: outdata = 32'd5708;
			59829: outdata = 32'd5707;
			59830: outdata = 32'd5706;
			59831: outdata = 32'd5705;
			59832: outdata = 32'd5704;
			59833: outdata = 32'd5703;
			59834: outdata = 32'd5702;
			59835: outdata = 32'd5701;
			59836: outdata = 32'd5700;
			59837: outdata = 32'd5699;
			59838: outdata = 32'd5698;
			59839: outdata = 32'd5697;
			59840: outdata = 32'd5696;
			59841: outdata = 32'd5695;
			59842: outdata = 32'd5694;
			59843: outdata = 32'd5693;
			59844: outdata = 32'd5692;
			59845: outdata = 32'd5691;
			59846: outdata = 32'd5690;
			59847: outdata = 32'd5689;
			59848: outdata = 32'd5688;
			59849: outdata = 32'd5687;
			59850: outdata = 32'd5686;
			59851: outdata = 32'd5685;
			59852: outdata = 32'd5684;
			59853: outdata = 32'd5683;
			59854: outdata = 32'd5682;
			59855: outdata = 32'd5681;
			59856: outdata = 32'd5680;
			59857: outdata = 32'd5679;
			59858: outdata = 32'd5678;
			59859: outdata = 32'd5677;
			59860: outdata = 32'd5676;
			59861: outdata = 32'd5675;
			59862: outdata = 32'd5674;
			59863: outdata = 32'd5673;
			59864: outdata = 32'd5672;
			59865: outdata = 32'd5671;
			59866: outdata = 32'd5670;
			59867: outdata = 32'd5669;
			59868: outdata = 32'd5668;
			59869: outdata = 32'd5667;
			59870: outdata = 32'd5666;
			59871: outdata = 32'd5665;
			59872: outdata = 32'd5664;
			59873: outdata = 32'd5663;
			59874: outdata = 32'd5662;
			59875: outdata = 32'd5661;
			59876: outdata = 32'd5660;
			59877: outdata = 32'd5659;
			59878: outdata = 32'd5658;
			59879: outdata = 32'd5657;
			59880: outdata = 32'd5656;
			59881: outdata = 32'd5655;
			59882: outdata = 32'd5654;
			59883: outdata = 32'd5653;
			59884: outdata = 32'd5652;
			59885: outdata = 32'd5651;
			59886: outdata = 32'd5650;
			59887: outdata = 32'd5649;
			59888: outdata = 32'd5648;
			59889: outdata = 32'd5647;
			59890: outdata = 32'd5646;
			59891: outdata = 32'd5645;
			59892: outdata = 32'd5644;
			59893: outdata = 32'd5643;
			59894: outdata = 32'd5642;
			59895: outdata = 32'd5641;
			59896: outdata = 32'd5640;
			59897: outdata = 32'd5639;
			59898: outdata = 32'd5638;
			59899: outdata = 32'd5637;
			59900: outdata = 32'd5636;
			59901: outdata = 32'd5635;
			59902: outdata = 32'd5634;
			59903: outdata = 32'd5633;
			59904: outdata = 32'd5632;
			59905: outdata = 32'd5631;
			59906: outdata = 32'd5630;
			59907: outdata = 32'd5629;
			59908: outdata = 32'd5628;
			59909: outdata = 32'd5627;
			59910: outdata = 32'd5626;
			59911: outdata = 32'd5625;
			59912: outdata = 32'd5624;
			59913: outdata = 32'd5623;
			59914: outdata = 32'd5622;
			59915: outdata = 32'd5621;
			59916: outdata = 32'd5620;
			59917: outdata = 32'd5619;
			59918: outdata = 32'd5618;
			59919: outdata = 32'd5617;
			59920: outdata = 32'd5616;
			59921: outdata = 32'd5615;
			59922: outdata = 32'd5614;
			59923: outdata = 32'd5613;
			59924: outdata = 32'd5612;
			59925: outdata = 32'd5611;
			59926: outdata = 32'd5610;
			59927: outdata = 32'd5609;
			59928: outdata = 32'd5608;
			59929: outdata = 32'd5607;
			59930: outdata = 32'd5606;
			59931: outdata = 32'd5605;
			59932: outdata = 32'd5604;
			59933: outdata = 32'd5603;
			59934: outdata = 32'd5602;
			59935: outdata = 32'd5601;
			59936: outdata = 32'd5600;
			59937: outdata = 32'd5599;
			59938: outdata = 32'd5598;
			59939: outdata = 32'd5597;
			59940: outdata = 32'd5596;
			59941: outdata = 32'd5595;
			59942: outdata = 32'd5594;
			59943: outdata = 32'd5593;
			59944: outdata = 32'd5592;
			59945: outdata = 32'd5591;
			59946: outdata = 32'd5590;
			59947: outdata = 32'd5589;
			59948: outdata = 32'd5588;
			59949: outdata = 32'd5587;
			59950: outdata = 32'd5586;
			59951: outdata = 32'd5585;
			59952: outdata = 32'd5584;
			59953: outdata = 32'd5583;
			59954: outdata = 32'd5582;
			59955: outdata = 32'd5581;
			59956: outdata = 32'd5580;
			59957: outdata = 32'd5579;
			59958: outdata = 32'd5578;
			59959: outdata = 32'd5577;
			59960: outdata = 32'd5576;
			59961: outdata = 32'd5575;
			59962: outdata = 32'd5574;
			59963: outdata = 32'd5573;
			59964: outdata = 32'd5572;
			59965: outdata = 32'd5571;
			59966: outdata = 32'd5570;
			59967: outdata = 32'd5569;
			59968: outdata = 32'd5568;
			59969: outdata = 32'd5567;
			59970: outdata = 32'd5566;
			59971: outdata = 32'd5565;
			59972: outdata = 32'd5564;
			59973: outdata = 32'd5563;
			59974: outdata = 32'd5562;
			59975: outdata = 32'd5561;
			59976: outdata = 32'd5560;
			59977: outdata = 32'd5559;
			59978: outdata = 32'd5558;
			59979: outdata = 32'd5557;
			59980: outdata = 32'd5556;
			59981: outdata = 32'd5555;
			59982: outdata = 32'd5554;
			59983: outdata = 32'd5553;
			59984: outdata = 32'd5552;
			59985: outdata = 32'd5551;
			59986: outdata = 32'd5550;
			59987: outdata = 32'd5549;
			59988: outdata = 32'd5548;
			59989: outdata = 32'd5547;
			59990: outdata = 32'd5546;
			59991: outdata = 32'd5545;
			59992: outdata = 32'd5544;
			59993: outdata = 32'd5543;
			59994: outdata = 32'd5542;
			59995: outdata = 32'd5541;
			59996: outdata = 32'd5540;
			59997: outdata = 32'd5539;
			59998: outdata = 32'd5538;
			59999: outdata = 32'd5537;
			60000: outdata = 32'd5536;
			60001: outdata = 32'd5535;
			60002: outdata = 32'd5534;
			60003: outdata = 32'd5533;
			60004: outdata = 32'd5532;
			60005: outdata = 32'd5531;
			60006: outdata = 32'd5530;
			60007: outdata = 32'd5529;
			60008: outdata = 32'd5528;
			60009: outdata = 32'd5527;
			60010: outdata = 32'd5526;
			60011: outdata = 32'd5525;
			60012: outdata = 32'd5524;
			60013: outdata = 32'd5523;
			60014: outdata = 32'd5522;
			60015: outdata = 32'd5521;
			60016: outdata = 32'd5520;
			60017: outdata = 32'd5519;
			60018: outdata = 32'd5518;
			60019: outdata = 32'd5517;
			60020: outdata = 32'd5516;
			60021: outdata = 32'd5515;
			60022: outdata = 32'd5514;
			60023: outdata = 32'd5513;
			60024: outdata = 32'd5512;
			60025: outdata = 32'd5511;
			60026: outdata = 32'd5510;
			60027: outdata = 32'd5509;
			60028: outdata = 32'd5508;
			60029: outdata = 32'd5507;
			60030: outdata = 32'd5506;
			60031: outdata = 32'd5505;
			60032: outdata = 32'd5504;
			60033: outdata = 32'd5503;
			60034: outdata = 32'd5502;
			60035: outdata = 32'd5501;
			60036: outdata = 32'd5500;
			60037: outdata = 32'd5499;
			60038: outdata = 32'd5498;
			60039: outdata = 32'd5497;
			60040: outdata = 32'd5496;
			60041: outdata = 32'd5495;
			60042: outdata = 32'd5494;
			60043: outdata = 32'd5493;
			60044: outdata = 32'd5492;
			60045: outdata = 32'd5491;
			60046: outdata = 32'd5490;
			60047: outdata = 32'd5489;
			60048: outdata = 32'd5488;
			60049: outdata = 32'd5487;
			60050: outdata = 32'd5486;
			60051: outdata = 32'd5485;
			60052: outdata = 32'd5484;
			60053: outdata = 32'd5483;
			60054: outdata = 32'd5482;
			60055: outdata = 32'd5481;
			60056: outdata = 32'd5480;
			60057: outdata = 32'd5479;
			60058: outdata = 32'd5478;
			60059: outdata = 32'd5477;
			60060: outdata = 32'd5476;
			60061: outdata = 32'd5475;
			60062: outdata = 32'd5474;
			60063: outdata = 32'd5473;
			60064: outdata = 32'd5472;
			60065: outdata = 32'd5471;
			60066: outdata = 32'd5470;
			60067: outdata = 32'd5469;
			60068: outdata = 32'd5468;
			60069: outdata = 32'd5467;
			60070: outdata = 32'd5466;
			60071: outdata = 32'd5465;
			60072: outdata = 32'd5464;
			60073: outdata = 32'd5463;
			60074: outdata = 32'd5462;
			60075: outdata = 32'd5461;
			60076: outdata = 32'd5460;
			60077: outdata = 32'd5459;
			60078: outdata = 32'd5458;
			60079: outdata = 32'd5457;
			60080: outdata = 32'd5456;
			60081: outdata = 32'd5455;
			60082: outdata = 32'd5454;
			60083: outdata = 32'd5453;
			60084: outdata = 32'd5452;
			60085: outdata = 32'd5451;
			60086: outdata = 32'd5450;
			60087: outdata = 32'd5449;
			60088: outdata = 32'd5448;
			60089: outdata = 32'd5447;
			60090: outdata = 32'd5446;
			60091: outdata = 32'd5445;
			60092: outdata = 32'd5444;
			60093: outdata = 32'd5443;
			60094: outdata = 32'd5442;
			60095: outdata = 32'd5441;
			60096: outdata = 32'd5440;
			60097: outdata = 32'd5439;
			60098: outdata = 32'd5438;
			60099: outdata = 32'd5437;
			60100: outdata = 32'd5436;
			60101: outdata = 32'd5435;
			60102: outdata = 32'd5434;
			60103: outdata = 32'd5433;
			60104: outdata = 32'd5432;
			60105: outdata = 32'd5431;
			60106: outdata = 32'd5430;
			60107: outdata = 32'd5429;
			60108: outdata = 32'd5428;
			60109: outdata = 32'd5427;
			60110: outdata = 32'd5426;
			60111: outdata = 32'd5425;
			60112: outdata = 32'd5424;
			60113: outdata = 32'd5423;
			60114: outdata = 32'd5422;
			60115: outdata = 32'd5421;
			60116: outdata = 32'd5420;
			60117: outdata = 32'd5419;
			60118: outdata = 32'd5418;
			60119: outdata = 32'd5417;
			60120: outdata = 32'd5416;
			60121: outdata = 32'd5415;
			60122: outdata = 32'd5414;
			60123: outdata = 32'd5413;
			60124: outdata = 32'd5412;
			60125: outdata = 32'd5411;
			60126: outdata = 32'd5410;
			60127: outdata = 32'd5409;
			60128: outdata = 32'd5408;
			60129: outdata = 32'd5407;
			60130: outdata = 32'd5406;
			60131: outdata = 32'd5405;
			60132: outdata = 32'd5404;
			60133: outdata = 32'd5403;
			60134: outdata = 32'd5402;
			60135: outdata = 32'd5401;
			60136: outdata = 32'd5400;
			60137: outdata = 32'd5399;
			60138: outdata = 32'd5398;
			60139: outdata = 32'd5397;
			60140: outdata = 32'd5396;
			60141: outdata = 32'd5395;
			60142: outdata = 32'd5394;
			60143: outdata = 32'd5393;
			60144: outdata = 32'd5392;
			60145: outdata = 32'd5391;
			60146: outdata = 32'd5390;
			60147: outdata = 32'd5389;
			60148: outdata = 32'd5388;
			60149: outdata = 32'd5387;
			60150: outdata = 32'd5386;
			60151: outdata = 32'd5385;
			60152: outdata = 32'd5384;
			60153: outdata = 32'd5383;
			60154: outdata = 32'd5382;
			60155: outdata = 32'd5381;
			60156: outdata = 32'd5380;
			60157: outdata = 32'd5379;
			60158: outdata = 32'd5378;
			60159: outdata = 32'd5377;
			60160: outdata = 32'd5376;
			60161: outdata = 32'd5375;
			60162: outdata = 32'd5374;
			60163: outdata = 32'd5373;
			60164: outdata = 32'd5372;
			60165: outdata = 32'd5371;
			60166: outdata = 32'd5370;
			60167: outdata = 32'd5369;
			60168: outdata = 32'd5368;
			60169: outdata = 32'd5367;
			60170: outdata = 32'd5366;
			60171: outdata = 32'd5365;
			60172: outdata = 32'd5364;
			60173: outdata = 32'd5363;
			60174: outdata = 32'd5362;
			60175: outdata = 32'd5361;
			60176: outdata = 32'd5360;
			60177: outdata = 32'd5359;
			60178: outdata = 32'd5358;
			60179: outdata = 32'd5357;
			60180: outdata = 32'd5356;
			60181: outdata = 32'd5355;
			60182: outdata = 32'd5354;
			60183: outdata = 32'd5353;
			60184: outdata = 32'd5352;
			60185: outdata = 32'd5351;
			60186: outdata = 32'd5350;
			60187: outdata = 32'd5349;
			60188: outdata = 32'd5348;
			60189: outdata = 32'd5347;
			60190: outdata = 32'd5346;
			60191: outdata = 32'd5345;
			60192: outdata = 32'd5344;
			60193: outdata = 32'd5343;
			60194: outdata = 32'd5342;
			60195: outdata = 32'd5341;
			60196: outdata = 32'd5340;
			60197: outdata = 32'd5339;
			60198: outdata = 32'd5338;
			60199: outdata = 32'd5337;
			60200: outdata = 32'd5336;
			60201: outdata = 32'd5335;
			60202: outdata = 32'd5334;
			60203: outdata = 32'd5333;
			60204: outdata = 32'd5332;
			60205: outdata = 32'd5331;
			60206: outdata = 32'd5330;
			60207: outdata = 32'd5329;
			60208: outdata = 32'd5328;
			60209: outdata = 32'd5327;
			60210: outdata = 32'd5326;
			60211: outdata = 32'd5325;
			60212: outdata = 32'd5324;
			60213: outdata = 32'd5323;
			60214: outdata = 32'd5322;
			60215: outdata = 32'd5321;
			60216: outdata = 32'd5320;
			60217: outdata = 32'd5319;
			60218: outdata = 32'd5318;
			60219: outdata = 32'd5317;
			60220: outdata = 32'd5316;
			60221: outdata = 32'd5315;
			60222: outdata = 32'd5314;
			60223: outdata = 32'd5313;
			60224: outdata = 32'd5312;
			60225: outdata = 32'd5311;
			60226: outdata = 32'd5310;
			60227: outdata = 32'd5309;
			60228: outdata = 32'd5308;
			60229: outdata = 32'd5307;
			60230: outdata = 32'd5306;
			60231: outdata = 32'd5305;
			60232: outdata = 32'd5304;
			60233: outdata = 32'd5303;
			60234: outdata = 32'd5302;
			60235: outdata = 32'd5301;
			60236: outdata = 32'd5300;
			60237: outdata = 32'd5299;
			60238: outdata = 32'd5298;
			60239: outdata = 32'd5297;
			60240: outdata = 32'd5296;
			60241: outdata = 32'd5295;
			60242: outdata = 32'd5294;
			60243: outdata = 32'd5293;
			60244: outdata = 32'd5292;
			60245: outdata = 32'd5291;
			60246: outdata = 32'd5290;
			60247: outdata = 32'd5289;
			60248: outdata = 32'd5288;
			60249: outdata = 32'd5287;
			60250: outdata = 32'd5286;
			60251: outdata = 32'd5285;
			60252: outdata = 32'd5284;
			60253: outdata = 32'd5283;
			60254: outdata = 32'd5282;
			60255: outdata = 32'd5281;
			60256: outdata = 32'd5280;
			60257: outdata = 32'd5279;
			60258: outdata = 32'd5278;
			60259: outdata = 32'd5277;
			60260: outdata = 32'd5276;
			60261: outdata = 32'd5275;
			60262: outdata = 32'd5274;
			60263: outdata = 32'd5273;
			60264: outdata = 32'd5272;
			60265: outdata = 32'd5271;
			60266: outdata = 32'd5270;
			60267: outdata = 32'd5269;
			60268: outdata = 32'd5268;
			60269: outdata = 32'd5267;
			60270: outdata = 32'd5266;
			60271: outdata = 32'd5265;
			60272: outdata = 32'd5264;
			60273: outdata = 32'd5263;
			60274: outdata = 32'd5262;
			60275: outdata = 32'd5261;
			60276: outdata = 32'd5260;
			60277: outdata = 32'd5259;
			60278: outdata = 32'd5258;
			60279: outdata = 32'd5257;
			60280: outdata = 32'd5256;
			60281: outdata = 32'd5255;
			60282: outdata = 32'd5254;
			60283: outdata = 32'd5253;
			60284: outdata = 32'd5252;
			60285: outdata = 32'd5251;
			60286: outdata = 32'd5250;
			60287: outdata = 32'd5249;
			60288: outdata = 32'd5248;
			60289: outdata = 32'd5247;
			60290: outdata = 32'd5246;
			60291: outdata = 32'd5245;
			60292: outdata = 32'd5244;
			60293: outdata = 32'd5243;
			60294: outdata = 32'd5242;
			60295: outdata = 32'd5241;
			60296: outdata = 32'd5240;
			60297: outdata = 32'd5239;
			60298: outdata = 32'd5238;
			60299: outdata = 32'd5237;
			60300: outdata = 32'd5236;
			60301: outdata = 32'd5235;
			60302: outdata = 32'd5234;
			60303: outdata = 32'd5233;
			60304: outdata = 32'd5232;
			60305: outdata = 32'd5231;
			60306: outdata = 32'd5230;
			60307: outdata = 32'd5229;
			60308: outdata = 32'd5228;
			60309: outdata = 32'd5227;
			60310: outdata = 32'd5226;
			60311: outdata = 32'd5225;
			60312: outdata = 32'd5224;
			60313: outdata = 32'd5223;
			60314: outdata = 32'd5222;
			60315: outdata = 32'd5221;
			60316: outdata = 32'd5220;
			60317: outdata = 32'd5219;
			60318: outdata = 32'd5218;
			60319: outdata = 32'd5217;
			60320: outdata = 32'd5216;
			60321: outdata = 32'd5215;
			60322: outdata = 32'd5214;
			60323: outdata = 32'd5213;
			60324: outdata = 32'd5212;
			60325: outdata = 32'd5211;
			60326: outdata = 32'd5210;
			60327: outdata = 32'd5209;
			60328: outdata = 32'd5208;
			60329: outdata = 32'd5207;
			60330: outdata = 32'd5206;
			60331: outdata = 32'd5205;
			60332: outdata = 32'd5204;
			60333: outdata = 32'd5203;
			60334: outdata = 32'd5202;
			60335: outdata = 32'd5201;
			60336: outdata = 32'd5200;
			60337: outdata = 32'd5199;
			60338: outdata = 32'd5198;
			60339: outdata = 32'd5197;
			60340: outdata = 32'd5196;
			60341: outdata = 32'd5195;
			60342: outdata = 32'd5194;
			60343: outdata = 32'd5193;
			60344: outdata = 32'd5192;
			60345: outdata = 32'd5191;
			60346: outdata = 32'd5190;
			60347: outdata = 32'd5189;
			60348: outdata = 32'd5188;
			60349: outdata = 32'd5187;
			60350: outdata = 32'd5186;
			60351: outdata = 32'd5185;
			60352: outdata = 32'd5184;
			60353: outdata = 32'd5183;
			60354: outdata = 32'd5182;
			60355: outdata = 32'd5181;
			60356: outdata = 32'd5180;
			60357: outdata = 32'd5179;
			60358: outdata = 32'd5178;
			60359: outdata = 32'd5177;
			60360: outdata = 32'd5176;
			60361: outdata = 32'd5175;
			60362: outdata = 32'd5174;
			60363: outdata = 32'd5173;
			60364: outdata = 32'd5172;
			60365: outdata = 32'd5171;
			60366: outdata = 32'd5170;
			60367: outdata = 32'd5169;
			60368: outdata = 32'd5168;
			60369: outdata = 32'd5167;
			60370: outdata = 32'd5166;
			60371: outdata = 32'd5165;
			60372: outdata = 32'd5164;
			60373: outdata = 32'd5163;
			60374: outdata = 32'd5162;
			60375: outdata = 32'd5161;
			60376: outdata = 32'd5160;
			60377: outdata = 32'd5159;
			60378: outdata = 32'd5158;
			60379: outdata = 32'd5157;
			60380: outdata = 32'd5156;
			60381: outdata = 32'd5155;
			60382: outdata = 32'd5154;
			60383: outdata = 32'd5153;
			60384: outdata = 32'd5152;
			60385: outdata = 32'd5151;
			60386: outdata = 32'd5150;
			60387: outdata = 32'd5149;
			60388: outdata = 32'd5148;
			60389: outdata = 32'd5147;
			60390: outdata = 32'd5146;
			60391: outdata = 32'd5145;
			60392: outdata = 32'd5144;
			60393: outdata = 32'd5143;
			60394: outdata = 32'd5142;
			60395: outdata = 32'd5141;
			60396: outdata = 32'd5140;
			60397: outdata = 32'd5139;
			60398: outdata = 32'd5138;
			60399: outdata = 32'd5137;
			60400: outdata = 32'd5136;
			60401: outdata = 32'd5135;
			60402: outdata = 32'd5134;
			60403: outdata = 32'd5133;
			60404: outdata = 32'd5132;
			60405: outdata = 32'd5131;
			60406: outdata = 32'd5130;
			60407: outdata = 32'd5129;
			60408: outdata = 32'd5128;
			60409: outdata = 32'd5127;
			60410: outdata = 32'd5126;
			60411: outdata = 32'd5125;
			60412: outdata = 32'd5124;
			60413: outdata = 32'd5123;
			60414: outdata = 32'd5122;
			60415: outdata = 32'd5121;
			60416: outdata = 32'd5120;
			60417: outdata = 32'd5119;
			60418: outdata = 32'd5118;
			60419: outdata = 32'd5117;
			60420: outdata = 32'd5116;
			60421: outdata = 32'd5115;
			60422: outdata = 32'd5114;
			60423: outdata = 32'd5113;
			60424: outdata = 32'd5112;
			60425: outdata = 32'd5111;
			60426: outdata = 32'd5110;
			60427: outdata = 32'd5109;
			60428: outdata = 32'd5108;
			60429: outdata = 32'd5107;
			60430: outdata = 32'd5106;
			60431: outdata = 32'd5105;
			60432: outdata = 32'd5104;
			60433: outdata = 32'd5103;
			60434: outdata = 32'd5102;
			60435: outdata = 32'd5101;
			60436: outdata = 32'd5100;
			60437: outdata = 32'd5099;
			60438: outdata = 32'd5098;
			60439: outdata = 32'd5097;
			60440: outdata = 32'd5096;
			60441: outdata = 32'd5095;
			60442: outdata = 32'd5094;
			60443: outdata = 32'd5093;
			60444: outdata = 32'd5092;
			60445: outdata = 32'd5091;
			60446: outdata = 32'd5090;
			60447: outdata = 32'd5089;
			60448: outdata = 32'd5088;
			60449: outdata = 32'd5087;
			60450: outdata = 32'd5086;
			60451: outdata = 32'd5085;
			60452: outdata = 32'd5084;
			60453: outdata = 32'd5083;
			60454: outdata = 32'd5082;
			60455: outdata = 32'd5081;
			60456: outdata = 32'd5080;
			60457: outdata = 32'd5079;
			60458: outdata = 32'd5078;
			60459: outdata = 32'd5077;
			60460: outdata = 32'd5076;
			60461: outdata = 32'd5075;
			60462: outdata = 32'd5074;
			60463: outdata = 32'd5073;
			60464: outdata = 32'd5072;
			60465: outdata = 32'd5071;
			60466: outdata = 32'd5070;
			60467: outdata = 32'd5069;
			60468: outdata = 32'd5068;
			60469: outdata = 32'd5067;
			60470: outdata = 32'd5066;
			60471: outdata = 32'd5065;
			60472: outdata = 32'd5064;
			60473: outdata = 32'd5063;
			60474: outdata = 32'd5062;
			60475: outdata = 32'd5061;
			60476: outdata = 32'd5060;
			60477: outdata = 32'd5059;
			60478: outdata = 32'd5058;
			60479: outdata = 32'd5057;
			60480: outdata = 32'd5056;
			60481: outdata = 32'd5055;
			60482: outdata = 32'd5054;
			60483: outdata = 32'd5053;
			60484: outdata = 32'd5052;
			60485: outdata = 32'd5051;
			60486: outdata = 32'd5050;
			60487: outdata = 32'd5049;
			60488: outdata = 32'd5048;
			60489: outdata = 32'd5047;
			60490: outdata = 32'd5046;
			60491: outdata = 32'd5045;
			60492: outdata = 32'd5044;
			60493: outdata = 32'd5043;
			60494: outdata = 32'd5042;
			60495: outdata = 32'd5041;
			60496: outdata = 32'd5040;
			60497: outdata = 32'd5039;
			60498: outdata = 32'd5038;
			60499: outdata = 32'd5037;
			60500: outdata = 32'd5036;
			60501: outdata = 32'd5035;
			60502: outdata = 32'd5034;
			60503: outdata = 32'd5033;
			60504: outdata = 32'd5032;
			60505: outdata = 32'd5031;
			60506: outdata = 32'd5030;
			60507: outdata = 32'd5029;
			60508: outdata = 32'd5028;
			60509: outdata = 32'd5027;
			60510: outdata = 32'd5026;
			60511: outdata = 32'd5025;
			60512: outdata = 32'd5024;
			60513: outdata = 32'd5023;
			60514: outdata = 32'd5022;
			60515: outdata = 32'd5021;
			60516: outdata = 32'd5020;
			60517: outdata = 32'd5019;
			60518: outdata = 32'd5018;
			60519: outdata = 32'd5017;
			60520: outdata = 32'd5016;
			60521: outdata = 32'd5015;
			60522: outdata = 32'd5014;
			60523: outdata = 32'd5013;
			60524: outdata = 32'd5012;
			60525: outdata = 32'd5011;
			60526: outdata = 32'd5010;
			60527: outdata = 32'd5009;
			60528: outdata = 32'd5008;
			60529: outdata = 32'd5007;
			60530: outdata = 32'd5006;
			60531: outdata = 32'd5005;
			60532: outdata = 32'd5004;
			60533: outdata = 32'd5003;
			60534: outdata = 32'd5002;
			60535: outdata = 32'd5001;
			60536: outdata = 32'd5000;
			60537: outdata = 32'd4999;
			60538: outdata = 32'd4998;
			60539: outdata = 32'd4997;
			60540: outdata = 32'd4996;
			60541: outdata = 32'd4995;
			60542: outdata = 32'd4994;
			60543: outdata = 32'd4993;
			60544: outdata = 32'd4992;
			60545: outdata = 32'd4991;
			60546: outdata = 32'd4990;
			60547: outdata = 32'd4989;
			60548: outdata = 32'd4988;
			60549: outdata = 32'd4987;
			60550: outdata = 32'd4986;
			60551: outdata = 32'd4985;
			60552: outdata = 32'd4984;
			60553: outdata = 32'd4983;
			60554: outdata = 32'd4982;
			60555: outdata = 32'd4981;
			60556: outdata = 32'd4980;
			60557: outdata = 32'd4979;
			60558: outdata = 32'd4978;
			60559: outdata = 32'd4977;
			60560: outdata = 32'd4976;
			60561: outdata = 32'd4975;
			60562: outdata = 32'd4974;
			60563: outdata = 32'd4973;
			60564: outdata = 32'd4972;
			60565: outdata = 32'd4971;
			60566: outdata = 32'd4970;
			60567: outdata = 32'd4969;
			60568: outdata = 32'd4968;
			60569: outdata = 32'd4967;
			60570: outdata = 32'd4966;
			60571: outdata = 32'd4965;
			60572: outdata = 32'd4964;
			60573: outdata = 32'd4963;
			60574: outdata = 32'd4962;
			60575: outdata = 32'd4961;
			60576: outdata = 32'd4960;
			60577: outdata = 32'd4959;
			60578: outdata = 32'd4958;
			60579: outdata = 32'd4957;
			60580: outdata = 32'd4956;
			60581: outdata = 32'd4955;
			60582: outdata = 32'd4954;
			60583: outdata = 32'd4953;
			60584: outdata = 32'd4952;
			60585: outdata = 32'd4951;
			60586: outdata = 32'd4950;
			60587: outdata = 32'd4949;
			60588: outdata = 32'd4948;
			60589: outdata = 32'd4947;
			60590: outdata = 32'd4946;
			60591: outdata = 32'd4945;
			60592: outdata = 32'd4944;
			60593: outdata = 32'd4943;
			60594: outdata = 32'd4942;
			60595: outdata = 32'd4941;
			60596: outdata = 32'd4940;
			60597: outdata = 32'd4939;
			60598: outdata = 32'd4938;
			60599: outdata = 32'd4937;
			60600: outdata = 32'd4936;
			60601: outdata = 32'd4935;
			60602: outdata = 32'd4934;
			60603: outdata = 32'd4933;
			60604: outdata = 32'd4932;
			60605: outdata = 32'd4931;
			60606: outdata = 32'd4930;
			60607: outdata = 32'd4929;
			60608: outdata = 32'd4928;
			60609: outdata = 32'd4927;
			60610: outdata = 32'd4926;
			60611: outdata = 32'd4925;
			60612: outdata = 32'd4924;
			60613: outdata = 32'd4923;
			60614: outdata = 32'd4922;
			60615: outdata = 32'd4921;
			60616: outdata = 32'd4920;
			60617: outdata = 32'd4919;
			60618: outdata = 32'd4918;
			60619: outdata = 32'd4917;
			60620: outdata = 32'd4916;
			60621: outdata = 32'd4915;
			60622: outdata = 32'd4914;
			60623: outdata = 32'd4913;
			60624: outdata = 32'd4912;
			60625: outdata = 32'd4911;
			60626: outdata = 32'd4910;
			60627: outdata = 32'd4909;
			60628: outdata = 32'd4908;
			60629: outdata = 32'd4907;
			60630: outdata = 32'd4906;
			60631: outdata = 32'd4905;
			60632: outdata = 32'd4904;
			60633: outdata = 32'd4903;
			60634: outdata = 32'd4902;
			60635: outdata = 32'd4901;
			60636: outdata = 32'd4900;
			60637: outdata = 32'd4899;
			60638: outdata = 32'd4898;
			60639: outdata = 32'd4897;
			60640: outdata = 32'd4896;
			60641: outdata = 32'd4895;
			60642: outdata = 32'd4894;
			60643: outdata = 32'd4893;
			60644: outdata = 32'd4892;
			60645: outdata = 32'd4891;
			60646: outdata = 32'd4890;
			60647: outdata = 32'd4889;
			60648: outdata = 32'd4888;
			60649: outdata = 32'd4887;
			60650: outdata = 32'd4886;
			60651: outdata = 32'd4885;
			60652: outdata = 32'd4884;
			60653: outdata = 32'd4883;
			60654: outdata = 32'd4882;
			60655: outdata = 32'd4881;
			60656: outdata = 32'd4880;
			60657: outdata = 32'd4879;
			60658: outdata = 32'd4878;
			60659: outdata = 32'd4877;
			60660: outdata = 32'd4876;
			60661: outdata = 32'd4875;
			60662: outdata = 32'd4874;
			60663: outdata = 32'd4873;
			60664: outdata = 32'd4872;
			60665: outdata = 32'd4871;
			60666: outdata = 32'd4870;
			60667: outdata = 32'd4869;
			60668: outdata = 32'd4868;
			60669: outdata = 32'd4867;
			60670: outdata = 32'd4866;
			60671: outdata = 32'd4865;
			60672: outdata = 32'd4864;
			60673: outdata = 32'd4863;
			60674: outdata = 32'd4862;
			60675: outdata = 32'd4861;
			60676: outdata = 32'd4860;
			60677: outdata = 32'd4859;
			60678: outdata = 32'd4858;
			60679: outdata = 32'd4857;
			60680: outdata = 32'd4856;
			60681: outdata = 32'd4855;
			60682: outdata = 32'd4854;
			60683: outdata = 32'd4853;
			60684: outdata = 32'd4852;
			60685: outdata = 32'd4851;
			60686: outdata = 32'd4850;
			60687: outdata = 32'd4849;
			60688: outdata = 32'd4848;
			60689: outdata = 32'd4847;
			60690: outdata = 32'd4846;
			60691: outdata = 32'd4845;
			60692: outdata = 32'd4844;
			60693: outdata = 32'd4843;
			60694: outdata = 32'd4842;
			60695: outdata = 32'd4841;
			60696: outdata = 32'd4840;
			60697: outdata = 32'd4839;
			60698: outdata = 32'd4838;
			60699: outdata = 32'd4837;
			60700: outdata = 32'd4836;
			60701: outdata = 32'd4835;
			60702: outdata = 32'd4834;
			60703: outdata = 32'd4833;
			60704: outdata = 32'd4832;
			60705: outdata = 32'd4831;
			60706: outdata = 32'd4830;
			60707: outdata = 32'd4829;
			60708: outdata = 32'd4828;
			60709: outdata = 32'd4827;
			60710: outdata = 32'd4826;
			60711: outdata = 32'd4825;
			60712: outdata = 32'd4824;
			60713: outdata = 32'd4823;
			60714: outdata = 32'd4822;
			60715: outdata = 32'd4821;
			60716: outdata = 32'd4820;
			60717: outdata = 32'd4819;
			60718: outdata = 32'd4818;
			60719: outdata = 32'd4817;
			60720: outdata = 32'd4816;
			60721: outdata = 32'd4815;
			60722: outdata = 32'd4814;
			60723: outdata = 32'd4813;
			60724: outdata = 32'd4812;
			60725: outdata = 32'd4811;
			60726: outdata = 32'd4810;
			60727: outdata = 32'd4809;
			60728: outdata = 32'd4808;
			60729: outdata = 32'd4807;
			60730: outdata = 32'd4806;
			60731: outdata = 32'd4805;
			60732: outdata = 32'd4804;
			60733: outdata = 32'd4803;
			60734: outdata = 32'd4802;
			60735: outdata = 32'd4801;
			60736: outdata = 32'd4800;
			60737: outdata = 32'd4799;
			60738: outdata = 32'd4798;
			60739: outdata = 32'd4797;
			60740: outdata = 32'd4796;
			60741: outdata = 32'd4795;
			60742: outdata = 32'd4794;
			60743: outdata = 32'd4793;
			60744: outdata = 32'd4792;
			60745: outdata = 32'd4791;
			60746: outdata = 32'd4790;
			60747: outdata = 32'd4789;
			60748: outdata = 32'd4788;
			60749: outdata = 32'd4787;
			60750: outdata = 32'd4786;
			60751: outdata = 32'd4785;
			60752: outdata = 32'd4784;
			60753: outdata = 32'd4783;
			60754: outdata = 32'd4782;
			60755: outdata = 32'd4781;
			60756: outdata = 32'd4780;
			60757: outdata = 32'd4779;
			60758: outdata = 32'd4778;
			60759: outdata = 32'd4777;
			60760: outdata = 32'd4776;
			60761: outdata = 32'd4775;
			60762: outdata = 32'd4774;
			60763: outdata = 32'd4773;
			60764: outdata = 32'd4772;
			60765: outdata = 32'd4771;
			60766: outdata = 32'd4770;
			60767: outdata = 32'd4769;
			60768: outdata = 32'd4768;
			60769: outdata = 32'd4767;
			60770: outdata = 32'd4766;
			60771: outdata = 32'd4765;
			60772: outdata = 32'd4764;
			60773: outdata = 32'd4763;
			60774: outdata = 32'd4762;
			60775: outdata = 32'd4761;
			60776: outdata = 32'd4760;
			60777: outdata = 32'd4759;
			60778: outdata = 32'd4758;
			60779: outdata = 32'd4757;
			60780: outdata = 32'd4756;
			60781: outdata = 32'd4755;
			60782: outdata = 32'd4754;
			60783: outdata = 32'd4753;
			60784: outdata = 32'd4752;
			60785: outdata = 32'd4751;
			60786: outdata = 32'd4750;
			60787: outdata = 32'd4749;
			60788: outdata = 32'd4748;
			60789: outdata = 32'd4747;
			60790: outdata = 32'd4746;
			60791: outdata = 32'd4745;
			60792: outdata = 32'd4744;
			60793: outdata = 32'd4743;
			60794: outdata = 32'd4742;
			60795: outdata = 32'd4741;
			60796: outdata = 32'd4740;
			60797: outdata = 32'd4739;
			60798: outdata = 32'd4738;
			60799: outdata = 32'd4737;
			60800: outdata = 32'd4736;
			60801: outdata = 32'd4735;
			60802: outdata = 32'd4734;
			60803: outdata = 32'd4733;
			60804: outdata = 32'd4732;
			60805: outdata = 32'd4731;
			60806: outdata = 32'd4730;
			60807: outdata = 32'd4729;
			60808: outdata = 32'd4728;
			60809: outdata = 32'd4727;
			60810: outdata = 32'd4726;
			60811: outdata = 32'd4725;
			60812: outdata = 32'd4724;
			60813: outdata = 32'd4723;
			60814: outdata = 32'd4722;
			60815: outdata = 32'd4721;
			60816: outdata = 32'd4720;
			60817: outdata = 32'd4719;
			60818: outdata = 32'd4718;
			60819: outdata = 32'd4717;
			60820: outdata = 32'd4716;
			60821: outdata = 32'd4715;
			60822: outdata = 32'd4714;
			60823: outdata = 32'd4713;
			60824: outdata = 32'd4712;
			60825: outdata = 32'd4711;
			60826: outdata = 32'd4710;
			60827: outdata = 32'd4709;
			60828: outdata = 32'd4708;
			60829: outdata = 32'd4707;
			60830: outdata = 32'd4706;
			60831: outdata = 32'd4705;
			60832: outdata = 32'd4704;
			60833: outdata = 32'd4703;
			60834: outdata = 32'd4702;
			60835: outdata = 32'd4701;
			60836: outdata = 32'd4700;
			60837: outdata = 32'd4699;
			60838: outdata = 32'd4698;
			60839: outdata = 32'd4697;
			60840: outdata = 32'd4696;
			60841: outdata = 32'd4695;
			60842: outdata = 32'd4694;
			60843: outdata = 32'd4693;
			60844: outdata = 32'd4692;
			60845: outdata = 32'd4691;
			60846: outdata = 32'd4690;
			60847: outdata = 32'd4689;
			60848: outdata = 32'd4688;
			60849: outdata = 32'd4687;
			60850: outdata = 32'd4686;
			60851: outdata = 32'd4685;
			60852: outdata = 32'd4684;
			60853: outdata = 32'd4683;
			60854: outdata = 32'd4682;
			60855: outdata = 32'd4681;
			60856: outdata = 32'd4680;
			60857: outdata = 32'd4679;
			60858: outdata = 32'd4678;
			60859: outdata = 32'd4677;
			60860: outdata = 32'd4676;
			60861: outdata = 32'd4675;
			60862: outdata = 32'd4674;
			60863: outdata = 32'd4673;
			60864: outdata = 32'd4672;
			60865: outdata = 32'd4671;
			60866: outdata = 32'd4670;
			60867: outdata = 32'd4669;
			60868: outdata = 32'd4668;
			60869: outdata = 32'd4667;
			60870: outdata = 32'd4666;
			60871: outdata = 32'd4665;
			60872: outdata = 32'd4664;
			60873: outdata = 32'd4663;
			60874: outdata = 32'd4662;
			60875: outdata = 32'd4661;
			60876: outdata = 32'd4660;
			60877: outdata = 32'd4659;
			60878: outdata = 32'd4658;
			60879: outdata = 32'd4657;
			60880: outdata = 32'd4656;
			60881: outdata = 32'd4655;
			60882: outdata = 32'd4654;
			60883: outdata = 32'd4653;
			60884: outdata = 32'd4652;
			60885: outdata = 32'd4651;
			60886: outdata = 32'd4650;
			60887: outdata = 32'd4649;
			60888: outdata = 32'd4648;
			60889: outdata = 32'd4647;
			60890: outdata = 32'd4646;
			60891: outdata = 32'd4645;
			60892: outdata = 32'd4644;
			60893: outdata = 32'd4643;
			60894: outdata = 32'd4642;
			60895: outdata = 32'd4641;
			60896: outdata = 32'd4640;
			60897: outdata = 32'd4639;
			60898: outdata = 32'd4638;
			60899: outdata = 32'd4637;
			60900: outdata = 32'd4636;
			60901: outdata = 32'd4635;
			60902: outdata = 32'd4634;
			60903: outdata = 32'd4633;
			60904: outdata = 32'd4632;
			60905: outdata = 32'd4631;
			60906: outdata = 32'd4630;
			60907: outdata = 32'd4629;
			60908: outdata = 32'd4628;
			60909: outdata = 32'd4627;
			60910: outdata = 32'd4626;
			60911: outdata = 32'd4625;
			60912: outdata = 32'd4624;
			60913: outdata = 32'd4623;
			60914: outdata = 32'd4622;
			60915: outdata = 32'd4621;
			60916: outdata = 32'd4620;
			60917: outdata = 32'd4619;
			60918: outdata = 32'd4618;
			60919: outdata = 32'd4617;
			60920: outdata = 32'd4616;
			60921: outdata = 32'd4615;
			60922: outdata = 32'd4614;
			60923: outdata = 32'd4613;
			60924: outdata = 32'd4612;
			60925: outdata = 32'd4611;
			60926: outdata = 32'd4610;
			60927: outdata = 32'd4609;
			60928: outdata = 32'd4608;
			60929: outdata = 32'd4607;
			60930: outdata = 32'd4606;
			60931: outdata = 32'd4605;
			60932: outdata = 32'd4604;
			60933: outdata = 32'd4603;
			60934: outdata = 32'd4602;
			60935: outdata = 32'd4601;
			60936: outdata = 32'd4600;
			60937: outdata = 32'd4599;
			60938: outdata = 32'd4598;
			60939: outdata = 32'd4597;
			60940: outdata = 32'd4596;
			60941: outdata = 32'd4595;
			60942: outdata = 32'd4594;
			60943: outdata = 32'd4593;
			60944: outdata = 32'd4592;
			60945: outdata = 32'd4591;
			60946: outdata = 32'd4590;
			60947: outdata = 32'd4589;
			60948: outdata = 32'd4588;
			60949: outdata = 32'd4587;
			60950: outdata = 32'd4586;
			60951: outdata = 32'd4585;
			60952: outdata = 32'd4584;
			60953: outdata = 32'd4583;
			60954: outdata = 32'd4582;
			60955: outdata = 32'd4581;
			60956: outdata = 32'd4580;
			60957: outdata = 32'd4579;
			60958: outdata = 32'd4578;
			60959: outdata = 32'd4577;
			60960: outdata = 32'd4576;
			60961: outdata = 32'd4575;
			60962: outdata = 32'd4574;
			60963: outdata = 32'd4573;
			60964: outdata = 32'd4572;
			60965: outdata = 32'd4571;
			60966: outdata = 32'd4570;
			60967: outdata = 32'd4569;
			60968: outdata = 32'd4568;
			60969: outdata = 32'd4567;
			60970: outdata = 32'd4566;
			60971: outdata = 32'd4565;
			60972: outdata = 32'd4564;
			60973: outdata = 32'd4563;
			60974: outdata = 32'd4562;
			60975: outdata = 32'd4561;
			60976: outdata = 32'd4560;
			60977: outdata = 32'd4559;
			60978: outdata = 32'd4558;
			60979: outdata = 32'd4557;
			60980: outdata = 32'd4556;
			60981: outdata = 32'd4555;
			60982: outdata = 32'd4554;
			60983: outdata = 32'd4553;
			60984: outdata = 32'd4552;
			60985: outdata = 32'd4551;
			60986: outdata = 32'd4550;
			60987: outdata = 32'd4549;
			60988: outdata = 32'd4548;
			60989: outdata = 32'd4547;
			60990: outdata = 32'd4546;
			60991: outdata = 32'd4545;
			60992: outdata = 32'd4544;
			60993: outdata = 32'd4543;
			60994: outdata = 32'd4542;
			60995: outdata = 32'd4541;
			60996: outdata = 32'd4540;
			60997: outdata = 32'd4539;
			60998: outdata = 32'd4538;
			60999: outdata = 32'd4537;
			61000: outdata = 32'd4536;
			61001: outdata = 32'd4535;
			61002: outdata = 32'd4534;
			61003: outdata = 32'd4533;
			61004: outdata = 32'd4532;
			61005: outdata = 32'd4531;
			61006: outdata = 32'd4530;
			61007: outdata = 32'd4529;
			61008: outdata = 32'd4528;
			61009: outdata = 32'd4527;
			61010: outdata = 32'd4526;
			61011: outdata = 32'd4525;
			61012: outdata = 32'd4524;
			61013: outdata = 32'd4523;
			61014: outdata = 32'd4522;
			61015: outdata = 32'd4521;
			61016: outdata = 32'd4520;
			61017: outdata = 32'd4519;
			61018: outdata = 32'd4518;
			61019: outdata = 32'd4517;
			61020: outdata = 32'd4516;
			61021: outdata = 32'd4515;
			61022: outdata = 32'd4514;
			61023: outdata = 32'd4513;
			61024: outdata = 32'd4512;
			61025: outdata = 32'd4511;
			61026: outdata = 32'd4510;
			61027: outdata = 32'd4509;
			61028: outdata = 32'd4508;
			61029: outdata = 32'd4507;
			61030: outdata = 32'd4506;
			61031: outdata = 32'd4505;
			61032: outdata = 32'd4504;
			61033: outdata = 32'd4503;
			61034: outdata = 32'd4502;
			61035: outdata = 32'd4501;
			61036: outdata = 32'd4500;
			61037: outdata = 32'd4499;
			61038: outdata = 32'd4498;
			61039: outdata = 32'd4497;
			61040: outdata = 32'd4496;
			61041: outdata = 32'd4495;
			61042: outdata = 32'd4494;
			61043: outdata = 32'd4493;
			61044: outdata = 32'd4492;
			61045: outdata = 32'd4491;
			61046: outdata = 32'd4490;
			61047: outdata = 32'd4489;
			61048: outdata = 32'd4488;
			61049: outdata = 32'd4487;
			61050: outdata = 32'd4486;
			61051: outdata = 32'd4485;
			61052: outdata = 32'd4484;
			61053: outdata = 32'd4483;
			61054: outdata = 32'd4482;
			61055: outdata = 32'd4481;
			61056: outdata = 32'd4480;
			61057: outdata = 32'd4479;
			61058: outdata = 32'd4478;
			61059: outdata = 32'd4477;
			61060: outdata = 32'd4476;
			61061: outdata = 32'd4475;
			61062: outdata = 32'd4474;
			61063: outdata = 32'd4473;
			61064: outdata = 32'd4472;
			61065: outdata = 32'd4471;
			61066: outdata = 32'd4470;
			61067: outdata = 32'd4469;
			61068: outdata = 32'd4468;
			61069: outdata = 32'd4467;
			61070: outdata = 32'd4466;
			61071: outdata = 32'd4465;
			61072: outdata = 32'd4464;
			61073: outdata = 32'd4463;
			61074: outdata = 32'd4462;
			61075: outdata = 32'd4461;
			61076: outdata = 32'd4460;
			61077: outdata = 32'd4459;
			61078: outdata = 32'd4458;
			61079: outdata = 32'd4457;
			61080: outdata = 32'd4456;
			61081: outdata = 32'd4455;
			61082: outdata = 32'd4454;
			61083: outdata = 32'd4453;
			61084: outdata = 32'd4452;
			61085: outdata = 32'd4451;
			61086: outdata = 32'd4450;
			61087: outdata = 32'd4449;
			61088: outdata = 32'd4448;
			61089: outdata = 32'd4447;
			61090: outdata = 32'd4446;
			61091: outdata = 32'd4445;
			61092: outdata = 32'd4444;
			61093: outdata = 32'd4443;
			61094: outdata = 32'd4442;
			61095: outdata = 32'd4441;
			61096: outdata = 32'd4440;
			61097: outdata = 32'd4439;
			61098: outdata = 32'd4438;
			61099: outdata = 32'd4437;
			61100: outdata = 32'd4436;
			61101: outdata = 32'd4435;
			61102: outdata = 32'd4434;
			61103: outdata = 32'd4433;
			61104: outdata = 32'd4432;
			61105: outdata = 32'd4431;
			61106: outdata = 32'd4430;
			61107: outdata = 32'd4429;
			61108: outdata = 32'd4428;
			61109: outdata = 32'd4427;
			61110: outdata = 32'd4426;
			61111: outdata = 32'd4425;
			61112: outdata = 32'd4424;
			61113: outdata = 32'd4423;
			61114: outdata = 32'd4422;
			61115: outdata = 32'd4421;
			61116: outdata = 32'd4420;
			61117: outdata = 32'd4419;
			61118: outdata = 32'd4418;
			61119: outdata = 32'd4417;
			61120: outdata = 32'd4416;
			61121: outdata = 32'd4415;
			61122: outdata = 32'd4414;
			61123: outdata = 32'd4413;
			61124: outdata = 32'd4412;
			61125: outdata = 32'd4411;
			61126: outdata = 32'd4410;
			61127: outdata = 32'd4409;
			61128: outdata = 32'd4408;
			61129: outdata = 32'd4407;
			61130: outdata = 32'd4406;
			61131: outdata = 32'd4405;
			61132: outdata = 32'd4404;
			61133: outdata = 32'd4403;
			61134: outdata = 32'd4402;
			61135: outdata = 32'd4401;
			61136: outdata = 32'd4400;
			61137: outdata = 32'd4399;
			61138: outdata = 32'd4398;
			61139: outdata = 32'd4397;
			61140: outdata = 32'd4396;
			61141: outdata = 32'd4395;
			61142: outdata = 32'd4394;
			61143: outdata = 32'd4393;
			61144: outdata = 32'd4392;
			61145: outdata = 32'd4391;
			61146: outdata = 32'd4390;
			61147: outdata = 32'd4389;
			61148: outdata = 32'd4388;
			61149: outdata = 32'd4387;
			61150: outdata = 32'd4386;
			61151: outdata = 32'd4385;
			61152: outdata = 32'd4384;
			61153: outdata = 32'd4383;
			61154: outdata = 32'd4382;
			61155: outdata = 32'd4381;
			61156: outdata = 32'd4380;
			61157: outdata = 32'd4379;
			61158: outdata = 32'd4378;
			61159: outdata = 32'd4377;
			61160: outdata = 32'd4376;
			61161: outdata = 32'd4375;
			61162: outdata = 32'd4374;
			61163: outdata = 32'd4373;
			61164: outdata = 32'd4372;
			61165: outdata = 32'd4371;
			61166: outdata = 32'd4370;
			61167: outdata = 32'd4369;
			61168: outdata = 32'd4368;
			61169: outdata = 32'd4367;
			61170: outdata = 32'd4366;
			61171: outdata = 32'd4365;
			61172: outdata = 32'd4364;
			61173: outdata = 32'd4363;
			61174: outdata = 32'd4362;
			61175: outdata = 32'd4361;
			61176: outdata = 32'd4360;
			61177: outdata = 32'd4359;
			61178: outdata = 32'd4358;
			61179: outdata = 32'd4357;
			61180: outdata = 32'd4356;
			61181: outdata = 32'd4355;
			61182: outdata = 32'd4354;
			61183: outdata = 32'd4353;
			61184: outdata = 32'd4352;
			61185: outdata = 32'd4351;
			61186: outdata = 32'd4350;
			61187: outdata = 32'd4349;
			61188: outdata = 32'd4348;
			61189: outdata = 32'd4347;
			61190: outdata = 32'd4346;
			61191: outdata = 32'd4345;
			61192: outdata = 32'd4344;
			61193: outdata = 32'd4343;
			61194: outdata = 32'd4342;
			61195: outdata = 32'd4341;
			61196: outdata = 32'd4340;
			61197: outdata = 32'd4339;
			61198: outdata = 32'd4338;
			61199: outdata = 32'd4337;
			61200: outdata = 32'd4336;
			61201: outdata = 32'd4335;
			61202: outdata = 32'd4334;
			61203: outdata = 32'd4333;
			61204: outdata = 32'd4332;
			61205: outdata = 32'd4331;
			61206: outdata = 32'd4330;
			61207: outdata = 32'd4329;
			61208: outdata = 32'd4328;
			61209: outdata = 32'd4327;
			61210: outdata = 32'd4326;
			61211: outdata = 32'd4325;
			61212: outdata = 32'd4324;
			61213: outdata = 32'd4323;
			61214: outdata = 32'd4322;
			61215: outdata = 32'd4321;
			61216: outdata = 32'd4320;
			61217: outdata = 32'd4319;
			61218: outdata = 32'd4318;
			61219: outdata = 32'd4317;
			61220: outdata = 32'd4316;
			61221: outdata = 32'd4315;
			61222: outdata = 32'd4314;
			61223: outdata = 32'd4313;
			61224: outdata = 32'd4312;
			61225: outdata = 32'd4311;
			61226: outdata = 32'd4310;
			61227: outdata = 32'd4309;
			61228: outdata = 32'd4308;
			61229: outdata = 32'd4307;
			61230: outdata = 32'd4306;
			61231: outdata = 32'd4305;
			61232: outdata = 32'd4304;
			61233: outdata = 32'd4303;
			61234: outdata = 32'd4302;
			61235: outdata = 32'd4301;
			61236: outdata = 32'd4300;
			61237: outdata = 32'd4299;
			61238: outdata = 32'd4298;
			61239: outdata = 32'd4297;
			61240: outdata = 32'd4296;
			61241: outdata = 32'd4295;
			61242: outdata = 32'd4294;
			61243: outdata = 32'd4293;
			61244: outdata = 32'd4292;
			61245: outdata = 32'd4291;
			61246: outdata = 32'd4290;
			61247: outdata = 32'd4289;
			61248: outdata = 32'd4288;
			61249: outdata = 32'd4287;
			61250: outdata = 32'd4286;
			61251: outdata = 32'd4285;
			61252: outdata = 32'd4284;
			61253: outdata = 32'd4283;
			61254: outdata = 32'd4282;
			61255: outdata = 32'd4281;
			61256: outdata = 32'd4280;
			61257: outdata = 32'd4279;
			61258: outdata = 32'd4278;
			61259: outdata = 32'd4277;
			61260: outdata = 32'd4276;
			61261: outdata = 32'd4275;
			61262: outdata = 32'd4274;
			61263: outdata = 32'd4273;
			61264: outdata = 32'd4272;
			61265: outdata = 32'd4271;
			61266: outdata = 32'd4270;
			61267: outdata = 32'd4269;
			61268: outdata = 32'd4268;
			61269: outdata = 32'd4267;
			61270: outdata = 32'd4266;
			61271: outdata = 32'd4265;
			61272: outdata = 32'd4264;
			61273: outdata = 32'd4263;
			61274: outdata = 32'd4262;
			61275: outdata = 32'd4261;
			61276: outdata = 32'd4260;
			61277: outdata = 32'd4259;
			61278: outdata = 32'd4258;
			61279: outdata = 32'd4257;
			61280: outdata = 32'd4256;
			61281: outdata = 32'd4255;
			61282: outdata = 32'd4254;
			61283: outdata = 32'd4253;
			61284: outdata = 32'd4252;
			61285: outdata = 32'd4251;
			61286: outdata = 32'd4250;
			61287: outdata = 32'd4249;
			61288: outdata = 32'd4248;
			61289: outdata = 32'd4247;
			61290: outdata = 32'd4246;
			61291: outdata = 32'd4245;
			61292: outdata = 32'd4244;
			61293: outdata = 32'd4243;
			61294: outdata = 32'd4242;
			61295: outdata = 32'd4241;
			61296: outdata = 32'd4240;
			61297: outdata = 32'd4239;
			61298: outdata = 32'd4238;
			61299: outdata = 32'd4237;
			61300: outdata = 32'd4236;
			61301: outdata = 32'd4235;
			61302: outdata = 32'd4234;
			61303: outdata = 32'd4233;
			61304: outdata = 32'd4232;
			61305: outdata = 32'd4231;
			61306: outdata = 32'd4230;
			61307: outdata = 32'd4229;
			61308: outdata = 32'd4228;
			61309: outdata = 32'd4227;
			61310: outdata = 32'd4226;
			61311: outdata = 32'd4225;
			61312: outdata = 32'd4224;
			61313: outdata = 32'd4223;
			61314: outdata = 32'd4222;
			61315: outdata = 32'd4221;
			61316: outdata = 32'd4220;
			61317: outdata = 32'd4219;
			61318: outdata = 32'd4218;
			61319: outdata = 32'd4217;
			61320: outdata = 32'd4216;
			61321: outdata = 32'd4215;
			61322: outdata = 32'd4214;
			61323: outdata = 32'd4213;
			61324: outdata = 32'd4212;
			61325: outdata = 32'd4211;
			61326: outdata = 32'd4210;
			61327: outdata = 32'd4209;
			61328: outdata = 32'd4208;
			61329: outdata = 32'd4207;
			61330: outdata = 32'd4206;
			61331: outdata = 32'd4205;
			61332: outdata = 32'd4204;
			61333: outdata = 32'd4203;
			61334: outdata = 32'd4202;
			61335: outdata = 32'd4201;
			61336: outdata = 32'd4200;
			61337: outdata = 32'd4199;
			61338: outdata = 32'd4198;
			61339: outdata = 32'd4197;
			61340: outdata = 32'd4196;
			61341: outdata = 32'd4195;
			61342: outdata = 32'd4194;
			61343: outdata = 32'd4193;
			61344: outdata = 32'd4192;
			61345: outdata = 32'd4191;
			61346: outdata = 32'd4190;
			61347: outdata = 32'd4189;
			61348: outdata = 32'd4188;
			61349: outdata = 32'd4187;
			61350: outdata = 32'd4186;
			61351: outdata = 32'd4185;
			61352: outdata = 32'd4184;
			61353: outdata = 32'd4183;
			61354: outdata = 32'd4182;
			61355: outdata = 32'd4181;
			61356: outdata = 32'd4180;
			61357: outdata = 32'd4179;
			61358: outdata = 32'd4178;
			61359: outdata = 32'd4177;
			61360: outdata = 32'd4176;
			61361: outdata = 32'd4175;
			61362: outdata = 32'd4174;
			61363: outdata = 32'd4173;
			61364: outdata = 32'd4172;
			61365: outdata = 32'd4171;
			61366: outdata = 32'd4170;
			61367: outdata = 32'd4169;
			61368: outdata = 32'd4168;
			61369: outdata = 32'd4167;
			61370: outdata = 32'd4166;
			61371: outdata = 32'd4165;
			61372: outdata = 32'd4164;
			61373: outdata = 32'd4163;
			61374: outdata = 32'd4162;
			61375: outdata = 32'd4161;
			61376: outdata = 32'd4160;
			61377: outdata = 32'd4159;
			61378: outdata = 32'd4158;
			61379: outdata = 32'd4157;
			61380: outdata = 32'd4156;
			61381: outdata = 32'd4155;
			61382: outdata = 32'd4154;
			61383: outdata = 32'd4153;
			61384: outdata = 32'd4152;
			61385: outdata = 32'd4151;
			61386: outdata = 32'd4150;
			61387: outdata = 32'd4149;
			61388: outdata = 32'd4148;
			61389: outdata = 32'd4147;
			61390: outdata = 32'd4146;
			61391: outdata = 32'd4145;
			61392: outdata = 32'd4144;
			61393: outdata = 32'd4143;
			61394: outdata = 32'd4142;
			61395: outdata = 32'd4141;
			61396: outdata = 32'd4140;
			61397: outdata = 32'd4139;
			61398: outdata = 32'd4138;
			61399: outdata = 32'd4137;
			61400: outdata = 32'd4136;
			61401: outdata = 32'd4135;
			61402: outdata = 32'd4134;
			61403: outdata = 32'd4133;
			61404: outdata = 32'd4132;
			61405: outdata = 32'd4131;
			61406: outdata = 32'd4130;
			61407: outdata = 32'd4129;
			61408: outdata = 32'd4128;
			61409: outdata = 32'd4127;
			61410: outdata = 32'd4126;
			61411: outdata = 32'd4125;
			61412: outdata = 32'd4124;
			61413: outdata = 32'd4123;
			61414: outdata = 32'd4122;
			61415: outdata = 32'd4121;
			61416: outdata = 32'd4120;
			61417: outdata = 32'd4119;
			61418: outdata = 32'd4118;
			61419: outdata = 32'd4117;
			61420: outdata = 32'd4116;
			61421: outdata = 32'd4115;
			61422: outdata = 32'd4114;
			61423: outdata = 32'd4113;
			61424: outdata = 32'd4112;
			61425: outdata = 32'd4111;
			61426: outdata = 32'd4110;
			61427: outdata = 32'd4109;
			61428: outdata = 32'd4108;
			61429: outdata = 32'd4107;
			61430: outdata = 32'd4106;
			61431: outdata = 32'd4105;
			61432: outdata = 32'd4104;
			61433: outdata = 32'd4103;
			61434: outdata = 32'd4102;
			61435: outdata = 32'd4101;
			61436: outdata = 32'd4100;
			61437: outdata = 32'd4099;
			61438: outdata = 32'd4098;
			61439: outdata = 32'd4097;
			61440: outdata = 32'd4096;
			61441: outdata = 32'd4095;
			61442: outdata = 32'd4094;
			61443: outdata = 32'd4093;
			61444: outdata = 32'd4092;
			61445: outdata = 32'd4091;
			61446: outdata = 32'd4090;
			61447: outdata = 32'd4089;
			61448: outdata = 32'd4088;
			61449: outdata = 32'd4087;
			61450: outdata = 32'd4086;
			61451: outdata = 32'd4085;
			61452: outdata = 32'd4084;
			61453: outdata = 32'd4083;
			61454: outdata = 32'd4082;
			61455: outdata = 32'd4081;
			61456: outdata = 32'd4080;
			61457: outdata = 32'd4079;
			61458: outdata = 32'd4078;
			61459: outdata = 32'd4077;
			61460: outdata = 32'd4076;
			61461: outdata = 32'd4075;
			61462: outdata = 32'd4074;
			61463: outdata = 32'd4073;
			61464: outdata = 32'd4072;
			61465: outdata = 32'd4071;
			61466: outdata = 32'd4070;
			61467: outdata = 32'd4069;
			61468: outdata = 32'd4068;
			61469: outdata = 32'd4067;
			61470: outdata = 32'd4066;
			61471: outdata = 32'd4065;
			61472: outdata = 32'd4064;
			61473: outdata = 32'd4063;
			61474: outdata = 32'd4062;
			61475: outdata = 32'd4061;
			61476: outdata = 32'd4060;
			61477: outdata = 32'd4059;
			61478: outdata = 32'd4058;
			61479: outdata = 32'd4057;
			61480: outdata = 32'd4056;
			61481: outdata = 32'd4055;
			61482: outdata = 32'd4054;
			61483: outdata = 32'd4053;
			61484: outdata = 32'd4052;
			61485: outdata = 32'd4051;
			61486: outdata = 32'd4050;
			61487: outdata = 32'd4049;
			61488: outdata = 32'd4048;
			61489: outdata = 32'd4047;
			61490: outdata = 32'd4046;
			61491: outdata = 32'd4045;
			61492: outdata = 32'd4044;
			61493: outdata = 32'd4043;
			61494: outdata = 32'd4042;
			61495: outdata = 32'd4041;
			61496: outdata = 32'd4040;
			61497: outdata = 32'd4039;
			61498: outdata = 32'd4038;
			61499: outdata = 32'd4037;
			61500: outdata = 32'd4036;
			61501: outdata = 32'd4035;
			61502: outdata = 32'd4034;
			61503: outdata = 32'd4033;
			61504: outdata = 32'd4032;
			61505: outdata = 32'd4031;
			61506: outdata = 32'd4030;
			61507: outdata = 32'd4029;
			61508: outdata = 32'd4028;
			61509: outdata = 32'd4027;
			61510: outdata = 32'd4026;
			61511: outdata = 32'd4025;
			61512: outdata = 32'd4024;
			61513: outdata = 32'd4023;
			61514: outdata = 32'd4022;
			61515: outdata = 32'd4021;
			61516: outdata = 32'd4020;
			61517: outdata = 32'd4019;
			61518: outdata = 32'd4018;
			61519: outdata = 32'd4017;
			61520: outdata = 32'd4016;
			61521: outdata = 32'd4015;
			61522: outdata = 32'd4014;
			61523: outdata = 32'd4013;
			61524: outdata = 32'd4012;
			61525: outdata = 32'd4011;
			61526: outdata = 32'd4010;
			61527: outdata = 32'd4009;
			61528: outdata = 32'd4008;
			61529: outdata = 32'd4007;
			61530: outdata = 32'd4006;
			61531: outdata = 32'd4005;
			61532: outdata = 32'd4004;
			61533: outdata = 32'd4003;
			61534: outdata = 32'd4002;
			61535: outdata = 32'd4001;
			61536: outdata = 32'd4000;
			61537: outdata = 32'd3999;
			61538: outdata = 32'd3998;
			61539: outdata = 32'd3997;
			61540: outdata = 32'd3996;
			61541: outdata = 32'd3995;
			61542: outdata = 32'd3994;
			61543: outdata = 32'd3993;
			61544: outdata = 32'd3992;
			61545: outdata = 32'd3991;
			61546: outdata = 32'd3990;
			61547: outdata = 32'd3989;
			61548: outdata = 32'd3988;
			61549: outdata = 32'd3987;
			61550: outdata = 32'd3986;
			61551: outdata = 32'd3985;
			61552: outdata = 32'd3984;
			61553: outdata = 32'd3983;
			61554: outdata = 32'd3982;
			61555: outdata = 32'd3981;
			61556: outdata = 32'd3980;
			61557: outdata = 32'd3979;
			61558: outdata = 32'd3978;
			61559: outdata = 32'd3977;
			61560: outdata = 32'd3976;
			61561: outdata = 32'd3975;
			61562: outdata = 32'd3974;
			61563: outdata = 32'd3973;
			61564: outdata = 32'd3972;
			61565: outdata = 32'd3971;
			61566: outdata = 32'd3970;
			61567: outdata = 32'd3969;
			61568: outdata = 32'd3968;
			61569: outdata = 32'd3967;
			61570: outdata = 32'd3966;
			61571: outdata = 32'd3965;
			61572: outdata = 32'd3964;
			61573: outdata = 32'd3963;
			61574: outdata = 32'd3962;
			61575: outdata = 32'd3961;
			61576: outdata = 32'd3960;
			61577: outdata = 32'd3959;
			61578: outdata = 32'd3958;
			61579: outdata = 32'd3957;
			61580: outdata = 32'd3956;
			61581: outdata = 32'd3955;
			61582: outdata = 32'd3954;
			61583: outdata = 32'd3953;
			61584: outdata = 32'd3952;
			61585: outdata = 32'd3951;
			61586: outdata = 32'd3950;
			61587: outdata = 32'd3949;
			61588: outdata = 32'd3948;
			61589: outdata = 32'd3947;
			61590: outdata = 32'd3946;
			61591: outdata = 32'd3945;
			61592: outdata = 32'd3944;
			61593: outdata = 32'd3943;
			61594: outdata = 32'd3942;
			61595: outdata = 32'd3941;
			61596: outdata = 32'd3940;
			61597: outdata = 32'd3939;
			61598: outdata = 32'd3938;
			61599: outdata = 32'd3937;
			61600: outdata = 32'd3936;
			61601: outdata = 32'd3935;
			61602: outdata = 32'd3934;
			61603: outdata = 32'd3933;
			61604: outdata = 32'd3932;
			61605: outdata = 32'd3931;
			61606: outdata = 32'd3930;
			61607: outdata = 32'd3929;
			61608: outdata = 32'd3928;
			61609: outdata = 32'd3927;
			61610: outdata = 32'd3926;
			61611: outdata = 32'd3925;
			61612: outdata = 32'd3924;
			61613: outdata = 32'd3923;
			61614: outdata = 32'd3922;
			61615: outdata = 32'd3921;
			61616: outdata = 32'd3920;
			61617: outdata = 32'd3919;
			61618: outdata = 32'd3918;
			61619: outdata = 32'd3917;
			61620: outdata = 32'd3916;
			61621: outdata = 32'd3915;
			61622: outdata = 32'd3914;
			61623: outdata = 32'd3913;
			61624: outdata = 32'd3912;
			61625: outdata = 32'd3911;
			61626: outdata = 32'd3910;
			61627: outdata = 32'd3909;
			61628: outdata = 32'd3908;
			61629: outdata = 32'd3907;
			61630: outdata = 32'd3906;
			61631: outdata = 32'd3905;
			61632: outdata = 32'd3904;
			61633: outdata = 32'd3903;
			61634: outdata = 32'd3902;
			61635: outdata = 32'd3901;
			61636: outdata = 32'd3900;
			61637: outdata = 32'd3899;
			61638: outdata = 32'd3898;
			61639: outdata = 32'd3897;
			61640: outdata = 32'd3896;
			61641: outdata = 32'd3895;
			61642: outdata = 32'd3894;
			61643: outdata = 32'd3893;
			61644: outdata = 32'd3892;
			61645: outdata = 32'd3891;
			61646: outdata = 32'd3890;
			61647: outdata = 32'd3889;
			61648: outdata = 32'd3888;
			61649: outdata = 32'd3887;
			61650: outdata = 32'd3886;
			61651: outdata = 32'd3885;
			61652: outdata = 32'd3884;
			61653: outdata = 32'd3883;
			61654: outdata = 32'd3882;
			61655: outdata = 32'd3881;
			61656: outdata = 32'd3880;
			61657: outdata = 32'd3879;
			61658: outdata = 32'd3878;
			61659: outdata = 32'd3877;
			61660: outdata = 32'd3876;
			61661: outdata = 32'd3875;
			61662: outdata = 32'd3874;
			61663: outdata = 32'd3873;
			61664: outdata = 32'd3872;
			61665: outdata = 32'd3871;
			61666: outdata = 32'd3870;
			61667: outdata = 32'd3869;
			61668: outdata = 32'd3868;
			61669: outdata = 32'd3867;
			61670: outdata = 32'd3866;
			61671: outdata = 32'd3865;
			61672: outdata = 32'd3864;
			61673: outdata = 32'd3863;
			61674: outdata = 32'd3862;
			61675: outdata = 32'd3861;
			61676: outdata = 32'd3860;
			61677: outdata = 32'd3859;
			61678: outdata = 32'd3858;
			61679: outdata = 32'd3857;
			61680: outdata = 32'd3856;
			61681: outdata = 32'd3855;
			61682: outdata = 32'd3854;
			61683: outdata = 32'd3853;
			61684: outdata = 32'd3852;
			61685: outdata = 32'd3851;
			61686: outdata = 32'd3850;
			61687: outdata = 32'd3849;
			61688: outdata = 32'd3848;
			61689: outdata = 32'd3847;
			61690: outdata = 32'd3846;
			61691: outdata = 32'd3845;
			61692: outdata = 32'd3844;
			61693: outdata = 32'd3843;
			61694: outdata = 32'd3842;
			61695: outdata = 32'd3841;
			61696: outdata = 32'd3840;
			61697: outdata = 32'd3839;
			61698: outdata = 32'd3838;
			61699: outdata = 32'd3837;
			61700: outdata = 32'd3836;
			61701: outdata = 32'd3835;
			61702: outdata = 32'd3834;
			61703: outdata = 32'd3833;
			61704: outdata = 32'd3832;
			61705: outdata = 32'd3831;
			61706: outdata = 32'd3830;
			61707: outdata = 32'd3829;
			61708: outdata = 32'd3828;
			61709: outdata = 32'd3827;
			61710: outdata = 32'd3826;
			61711: outdata = 32'd3825;
			61712: outdata = 32'd3824;
			61713: outdata = 32'd3823;
			61714: outdata = 32'd3822;
			61715: outdata = 32'd3821;
			61716: outdata = 32'd3820;
			61717: outdata = 32'd3819;
			61718: outdata = 32'd3818;
			61719: outdata = 32'd3817;
			61720: outdata = 32'd3816;
			61721: outdata = 32'd3815;
			61722: outdata = 32'd3814;
			61723: outdata = 32'd3813;
			61724: outdata = 32'd3812;
			61725: outdata = 32'd3811;
			61726: outdata = 32'd3810;
			61727: outdata = 32'd3809;
			61728: outdata = 32'd3808;
			61729: outdata = 32'd3807;
			61730: outdata = 32'd3806;
			61731: outdata = 32'd3805;
			61732: outdata = 32'd3804;
			61733: outdata = 32'd3803;
			61734: outdata = 32'd3802;
			61735: outdata = 32'd3801;
			61736: outdata = 32'd3800;
			61737: outdata = 32'd3799;
			61738: outdata = 32'd3798;
			61739: outdata = 32'd3797;
			61740: outdata = 32'd3796;
			61741: outdata = 32'd3795;
			61742: outdata = 32'd3794;
			61743: outdata = 32'd3793;
			61744: outdata = 32'd3792;
			61745: outdata = 32'd3791;
			61746: outdata = 32'd3790;
			61747: outdata = 32'd3789;
			61748: outdata = 32'd3788;
			61749: outdata = 32'd3787;
			61750: outdata = 32'd3786;
			61751: outdata = 32'd3785;
			61752: outdata = 32'd3784;
			61753: outdata = 32'd3783;
			61754: outdata = 32'd3782;
			61755: outdata = 32'd3781;
			61756: outdata = 32'd3780;
			61757: outdata = 32'd3779;
			61758: outdata = 32'd3778;
			61759: outdata = 32'd3777;
			61760: outdata = 32'd3776;
			61761: outdata = 32'd3775;
			61762: outdata = 32'd3774;
			61763: outdata = 32'd3773;
			61764: outdata = 32'd3772;
			61765: outdata = 32'd3771;
			61766: outdata = 32'd3770;
			61767: outdata = 32'd3769;
			61768: outdata = 32'd3768;
			61769: outdata = 32'd3767;
			61770: outdata = 32'd3766;
			61771: outdata = 32'd3765;
			61772: outdata = 32'd3764;
			61773: outdata = 32'd3763;
			61774: outdata = 32'd3762;
			61775: outdata = 32'd3761;
			61776: outdata = 32'd3760;
			61777: outdata = 32'd3759;
			61778: outdata = 32'd3758;
			61779: outdata = 32'd3757;
			61780: outdata = 32'd3756;
			61781: outdata = 32'd3755;
			61782: outdata = 32'd3754;
			61783: outdata = 32'd3753;
			61784: outdata = 32'd3752;
			61785: outdata = 32'd3751;
			61786: outdata = 32'd3750;
			61787: outdata = 32'd3749;
			61788: outdata = 32'd3748;
			61789: outdata = 32'd3747;
			61790: outdata = 32'd3746;
			61791: outdata = 32'd3745;
			61792: outdata = 32'd3744;
			61793: outdata = 32'd3743;
			61794: outdata = 32'd3742;
			61795: outdata = 32'd3741;
			61796: outdata = 32'd3740;
			61797: outdata = 32'd3739;
			61798: outdata = 32'd3738;
			61799: outdata = 32'd3737;
			61800: outdata = 32'd3736;
			61801: outdata = 32'd3735;
			61802: outdata = 32'd3734;
			61803: outdata = 32'd3733;
			61804: outdata = 32'd3732;
			61805: outdata = 32'd3731;
			61806: outdata = 32'd3730;
			61807: outdata = 32'd3729;
			61808: outdata = 32'd3728;
			61809: outdata = 32'd3727;
			61810: outdata = 32'd3726;
			61811: outdata = 32'd3725;
			61812: outdata = 32'd3724;
			61813: outdata = 32'd3723;
			61814: outdata = 32'd3722;
			61815: outdata = 32'd3721;
			61816: outdata = 32'd3720;
			61817: outdata = 32'd3719;
			61818: outdata = 32'd3718;
			61819: outdata = 32'd3717;
			61820: outdata = 32'd3716;
			61821: outdata = 32'd3715;
			61822: outdata = 32'd3714;
			61823: outdata = 32'd3713;
			61824: outdata = 32'd3712;
			61825: outdata = 32'd3711;
			61826: outdata = 32'd3710;
			61827: outdata = 32'd3709;
			61828: outdata = 32'd3708;
			61829: outdata = 32'd3707;
			61830: outdata = 32'd3706;
			61831: outdata = 32'd3705;
			61832: outdata = 32'd3704;
			61833: outdata = 32'd3703;
			61834: outdata = 32'd3702;
			61835: outdata = 32'd3701;
			61836: outdata = 32'd3700;
			61837: outdata = 32'd3699;
			61838: outdata = 32'd3698;
			61839: outdata = 32'd3697;
			61840: outdata = 32'd3696;
			61841: outdata = 32'd3695;
			61842: outdata = 32'd3694;
			61843: outdata = 32'd3693;
			61844: outdata = 32'd3692;
			61845: outdata = 32'd3691;
			61846: outdata = 32'd3690;
			61847: outdata = 32'd3689;
			61848: outdata = 32'd3688;
			61849: outdata = 32'd3687;
			61850: outdata = 32'd3686;
			61851: outdata = 32'd3685;
			61852: outdata = 32'd3684;
			61853: outdata = 32'd3683;
			61854: outdata = 32'd3682;
			61855: outdata = 32'd3681;
			61856: outdata = 32'd3680;
			61857: outdata = 32'd3679;
			61858: outdata = 32'd3678;
			61859: outdata = 32'd3677;
			61860: outdata = 32'd3676;
			61861: outdata = 32'd3675;
			61862: outdata = 32'd3674;
			61863: outdata = 32'd3673;
			61864: outdata = 32'd3672;
			61865: outdata = 32'd3671;
			61866: outdata = 32'd3670;
			61867: outdata = 32'd3669;
			61868: outdata = 32'd3668;
			61869: outdata = 32'd3667;
			61870: outdata = 32'd3666;
			61871: outdata = 32'd3665;
			61872: outdata = 32'd3664;
			61873: outdata = 32'd3663;
			61874: outdata = 32'd3662;
			61875: outdata = 32'd3661;
			61876: outdata = 32'd3660;
			61877: outdata = 32'd3659;
			61878: outdata = 32'd3658;
			61879: outdata = 32'd3657;
			61880: outdata = 32'd3656;
			61881: outdata = 32'd3655;
			61882: outdata = 32'd3654;
			61883: outdata = 32'd3653;
			61884: outdata = 32'd3652;
			61885: outdata = 32'd3651;
			61886: outdata = 32'd3650;
			61887: outdata = 32'd3649;
			61888: outdata = 32'd3648;
			61889: outdata = 32'd3647;
			61890: outdata = 32'd3646;
			61891: outdata = 32'd3645;
			61892: outdata = 32'd3644;
			61893: outdata = 32'd3643;
			61894: outdata = 32'd3642;
			61895: outdata = 32'd3641;
			61896: outdata = 32'd3640;
			61897: outdata = 32'd3639;
			61898: outdata = 32'd3638;
			61899: outdata = 32'd3637;
			61900: outdata = 32'd3636;
			61901: outdata = 32'd3635;
			61902: outdata = 32'd3634;
			61903: outdata = 32'd3633;
			61904: outdata = 32'd3632;
			61905: outdata = 32'd3631;
			61906: outdata = 32'd3630;
			61907: outdata = 32'd3629;
			61908: outdata = 32'd3628;
			61909: outdata = 32'd3627;
			61910: outdata = 32'd3626;
			61911: outdata = 32'd3625;
			61912: outdata = 32'd3624;
			61913: outdata = 32'd3623;
			61914: outdata = 32'd3622;
			61915: outdata = 32'd3621;
			61916: outdata = 32'd3620;
			61917: outdata = 32'd3619;
			61918: outdata = 32'd3618;
			61919: outdata = 32'd3617;
			61920: outdata = 32'd3616;
			61921: outdata = 32'd3615;
			61922: outdata = 32'd3614;
			61923: outdata = 32'd3613;
			61924: outdata = 32'd3612;
			61925: outdata = 32'd3611;
			61926: outdata = 32'd3610;
			61927: outdata = 32'd3609;
			61928: outdata = 32'd3608;
			61929: outdata = 32'd3607;
			61930: outdata = 32'd3606;
			61931: outdata = 32'd3605;
			61932: outdata = 32'd3604;
			61933: outdata = 32'd3603;
			61934: outdata = 32'd3602;
			61935: outdata = 32'd3601;
			61936: outdata = 32'd3600;
			61937: outdata = 32'd3599;
			61938: outdata = 32'd3598;
			61939: outdata = 32'd3597;
			61940: outdata = 32'd3596;
			61941: outdata = 32'd3595;
			61942: outdata = 32'd3594;
			61943: outdata = 32'd3593;
			61944: outdata = 32'd3592;
			61945: outdata = 32'd3591;
			61946: outdata = 32'd3590;
			61947: outdata = 32'd3589;
			61948: outdata = 32'd3588;
			61949: outdata = 32'd3587;
			61950: outdata = 32'd3586;
			61951: outdata = 32'd3585;
			61952: outdata = 32'd3584;
			61953: outdata = 32'd3583;
			61954: outdata = 32'd3582;
			61955: outdata = 32'd3581;
			61956: outdata = 32'd3580;
			61957: outdata = 32'd3579;
			61958: outdata = 32'd3578;
			61959: outdata = 32'd3577;
			61960: outdata = 32'd3576;
			61961: outdata = 32'd3575;
			61962: outdata = 32'd3574;
			61963: outdata = 32'd3573;
			61964: outdata = 32'd3572;
			61965: outdata = 32'd3571;
			61966: outdata = 32'd3570;
			61967: outdata = 32'd3569;
			61968: outdata = 32'd3568;
			61969: outdata = 32'd3567;
			61970: outdata = 32'd3566;
			61971: outdata = 32'd3565;
			61972: outdata = 32'd3564;
			61973: outdata = 32'd3563;
			61974: outdata = 32'd3562;
			61975: outdata = 32'd3561;
			61976: outdata = 32'd3560;
			61977: outdata = 32'd3559;
			61978: outdata = 32'd3558;
			61979: outdata = 32'd3557;
			61980: outdata = 32'd3556;
			61981: outdata = 32'd3555;
			61982: outdata = 32'd3554;
			61983: outdata = 32'd3553;
			61984: outdata = 32'd3552;
			61985: outdata = 32'd3551;
			61986: outdata = 32'd3550;
			61987: outdata = 32'd3549;
			61988: outdata = 32'd3548;
			61989: outdata = 32'd3547;
			61990: outdata = 32'd3546;
			61991: outdata = 32'd3545;
			61992: outdata = 32'd3544;
			61993: outdata = 32'd3543;
			61994: outdata = 32'd3542;
			61995: outdata = 32'd3541;
			61996: outdata = 32'd3540;
			61997: outdata = 32'd3539;
			61998: outdata = 32'd3538;
			61999: outdata = 32'd3537;
			62000: outdata = 32'd3536;
			62001: outdata = 32'd3535;
			62002: outdata = 32'd3534;
			62003: outdata = 32'd3533;
			62004: outdata = 32'd3532;
			62005: outdata = 32'd3531;
			62006: outdata = 32'd3530;
			62007: outdata = 32'd3529;
			62008: outdata = 32'd3528;
			62009: outdata = 32'd3527;
			62010: outdata = 32'd3526;
			62011: outdata = 32'd3525;
			62012: outdata = 32'd3524;
			62013: outdata = 32'd3523;
			62014: outdata = 32'd3522;
			62015: outdata = 32'd3521;
			62016: outdata = 32'd3520;
			62017: outdata = 32'd3519;
			62018: outdata = 32'd3518;
			62019: outdata = 32'd3517;
			62020: outdata = 32'd3516;
			62021: outdata = 32'd3515;
			62022: outdata = 32'd3514;
			62023: outdata = 32'd3513;
			62024: outdata = 32'd3512;
			62025: outdata = 32'd3511;
			62026: outdata = 32'd3510;
			62027: outdata = 32'd3509;
			62028: outdata = 32'd3508;
			62029: outdata = 32'd3507;
			62030: outdata = 32'd3506;
			62031: outdata = 32'd3505;
			62032: outdata = 32'd3504;
			62033: outdata = 32'd3503;
			62034: outdata = 32'd3502;
			62035: outdata = 32'd3501;
			62036: outdata = 32'd3500;
			62037: outdata = 32'd3499;
			62038: outdata = 32'd3498;
			62039: outdata = 32'd3497;
			62040: outdata = 32'd3496;
			62041: outdata = 32'd3495;
			62042: outdata = 32'd3494;
			62043: outdata = 32'd3493;
			62044: outdata = 32'd3492;
			62045: outdata = 32'd3491;
			62046: outdata = 32'd3490;
			62047: outdata = 32'd3489;
			62048: outdata = 32'd3488;
			62049: outdata = 32'd3487;
			62050: outdata = 32'd3486;
			62051: outdata = 32'd3485;
			62052: outdata = 32'd3484;
			62053: outdata = 32'd3483;
			62054: outdata = 32'd3482;
			62055: outdata = 32'd3481;
			62056: outdata = 32'd3480;
			62057: outdata = 32'd3479;
			62058: outdata = 32'd3478;
			62059: outdata = 32'd3477;
			62060: outdata = 32'd3476;
			62061: outdata = 32'd3475;
			62062: outdata = 32'd3474;
			62063: outdata = 32'd3473;
			62064: outdata = 32'd3472;
			62065: outdata = 32'd3471;
			62066: outdata = 32'd3470;
			62067: outdata = 32'd3469;
			62068: outdata = 32'd3468;
			62069: outdata = 32'd3467;
			62070: outdata = 32'd3466;
			62071: outdata = 32'd3465;
			62072: outdata = 32'd3464;
			62073: outdata = 32'd3463;
			62074: outdata = 32'd3462;
			62075: outdata = 32'd3461;
			62076: outdata = 32'd3460;
			62077: outdata = 32'd3459;
			62078: outdata = 32'd3458;
			62079: outdata = 32'd3457;
			62080: outdata = 32'd3456;
			62081: outdata = 32'd3455;
			62082: outdata = 32'd3454;
			62083: outdata = 32'd3453;
			62084: outdata = 32'd3452;
			62085: outdata = 32'd3451;
			62086: outdata = 32'd3450;
			62087: outdata = 32'd3449;
			62088: outdata = 32'd3448;
			62089: outdata = 32'd3447;
			62090: outdata = 32'd3446;
			62091: outdata = 32'd3445;
			62092: outdata = 32'd3444;
			62093: outdata = 32'd3443;
			62094: outdata = 32'd3442;
			62095: outdata = 32'd3441;
			62096: outdata = 32'd3440;
			62097: outdata = 32'd3439;
			62098: outdata = 32'd3438;
			62099: outdata = 32'd3437;
			62100: outdata = 32'd3436;
			62101: outdata = 32'd3435;
			62102: outdata = 32'd3434;
			62103: outdata = 32'd3433;
			62104: outdata = 32'd3432;
			62105: outdata = 32'd3431;
			62106: outdata = 32'd3430;
			62107: outdata = 32'd3429;
			62108: outdata = 32'd3428;
			62109: outdata = 32'd3427;
			62110: outdata = 32'd3426;
			62111: outdata = 32'd3425;
			62112: outdata = 32'd3424;
			62113: outdata = 32'd3423;
			62114: outdata = 32'd3422;
			62115: outdata = 32'd3421;
			62116: outdata = 32'd3420;
			62117: outdata = 32'd3419;
			62118: outdata = 32'd3418;
			62119: outdata = 32'd3417;
			62120: outdata = 32'd3416;
			62121: outdata = 32'd3415;
			62122: outdata = 32'd3414;
			62123: outdata = 32'd3413;
			62124: outdata = 32'd3412;
			62125: outdata = 32'd3411;
			62126: outdata = 32'd3410;
			62127: outdata = 32'd3409;
			62128: outdata = 32'd3408;
			62129: outdata = 32'd3407;
			62130: outdata = 32'd3406;
			62131: outdata = 32'd3405;
			62132: outdata = 32'd3404;
			62133: outdata = 32'd3403;
			62134: outdata = 32'd3402;
			62135: outdata = 32'd3401;
			62136: outdata = 32'd3400;
			62137: outdata = 32'd3399;
			62138: outdata = 32'd3398;
			62139: outdata = 32'd3397;
			62140: outdata = 32'd3396;
			62141: outdata = 32'd3395;
			62142: outdata = 32'd3394;
			62143: outdata = 32'd3393;
			62144: outdata = 32'd3392;
			62145: outdata = 32'd3391;
			62146: outdata = 32'd3390;
			62147: outdata = 32'd3389;
			62148: outdata = 32'd3388;
			62149: outdata = 32'd3387;
			62150: outdata = 32'd3386;
			62151: outdata = 32'd3385;
			62152: outdata = 32'd3384;
			62153: outdata = 32'd3383;
			62154: outdata = 32'd3382;
			62155: outdata = 32'd3381;
			62156: outdata = 32'd3380;
			62157: outdata = 32'd3379;
			62158: outdata = 32'd3378;
			62159: outdata = 32'd3377;
			62160: outdata = 32'd3376;
			62161: outdata = 32'd3375;
			62162: outdata = 32'd3374;
			62163: outdata = 32'd3373;
			62164: outdata = 32'd3372;
			62165: outdata = 32'd3371;
			62166: outdata = 32'd3370;
			62167: outdata = 32'd3369;
			62168: outdata = 32'd3368;
			62169: outdata = 32'd3367;
			62170: outdata = 32'd3366;
			62171: outdata = 32'd3365;
			62172: outdata = 32'd3364;
			62173: outdata = 32'd3363;
			62174: outdata = 32'd3362;
			62175: outdata = 32'd3361;
			62176: outdata = 32'd3360;
			62177: outdata = 32'd3359;
			62178: outdata = 32'd3358;
			62179: outdata = 32'd3357;
			62180: outdata = 32'd3356;
			62181: outdata = 32'd3355;
			62182: outdata = 32'd3354;
			62183: outdata = 32'd3353;
			62184: outdata = 32'd3352;
			62185: outdata = 32'd3351;
			62186: outdata = 32'd3350;
			62187: outdata = 32'd3349;
			62188: outdata = 32'd3348;
			62189: outdata = 32'd3347;
			62190: outdata = 32'd3346;
			62191: outdata = 32'd3345;
			62192: outdata = 32'd3344;
			62193: outdata = 32'd3343;
			62194: outdata = 32'd3342;
			62195: outdata = 32'd3341;
			62196: outdata = 32'd3340;
			62197: outdata = 32'd3339;
			62198: outdata = 32'd3338;
			62199: outdata = 32'd3337;
			62200: outdata = 32'd3336;
			62201: outdata = 32'd3335;
			62202: outdata = 32'd3334;
			62203: outdata = 32'd3333;
			62204: outdata = 32'd3332;
			62205: outdata = 32'd3331;
			62206: outdata = 32'd3330;
			62207: outdata = 32'd3329;
			62208: outdata = 32'd3328;
			62209: outdata = 32'd3327;
			62210: outdata = 32'd3326;
			62211: outdata = 32'd3325;
			62212: outdata = 32'd3324;
			62213: outdata = 32'd3323;
			62214: outdata = 32'd3322;
			62215: outdata = 32'd3321;
			62216: outdata = 32'd3320;
			62217: outdata = 32'd3319;
			62218: outdata = 32'd3318;
			62219: outdata = 32'd3317;
			62220: outdata = 32'd3316;
			62221: outdata = 32'd3315;
			62222: outdata = 32'd3314;
			62223: outdata = 32'd3313;
			62224: outdata = 32'd3312;
			62225: outdata = 32'd3311;
			62226: outdata = 32'd3310;
			62227: outdata = 32'd3309;
			62228: outdata = 32'd3308;
			62229: outdata = 32'd3307;
			62230: outdata = 32'd3306;
			62231: outdata = 32'd3305;
			62232: outdata = 32'd3304;
			62233: outdata = 32'd3303;
			62234: outdata = 32'd3302;
			62235: outdata = 32'd3301;
			62236: outdata = 32'd3300;
			62237: outdata = 32'd3299;
			62238: outdata = 32'd3298;
			62239: outdata = 32'd3297;
			62240: outdata = 32'd3296;
			62241: outdata = 32'd3295;
			62242: outdata = 32'd3294;
			62243: outdata = 32'd3293;
			62244: outdata = 32'd3292;
			62245: outdata = 32'd3291;
			62246: outdata = 32'd3290;
			62247: outdata = 32'd3289;
			62248: outdata = 32'd3288;
			62249: outdata = 32'd3287;
			62250: outdata = 32'd3286;
			62251: outdata = 32'd3285;
			62252: outdata = 32'd3284;
			62253: outdata = 32'd3283;
			62254: outdata = 32'd3282;
			62255: outdata = 32'd3281;
			62256: outdata = 32'd3280;
			62257: outdata = 32'd3279;
			62258: outdata = 32'd3278;
			62259: outdata = 32'd3277;
			62260: outdata = 32'd3276;
			62261: outdata = 32'd3275;
			62262: outdata = 32'd3274;
			62263: outdata = 32'd3273;
			62264: outdata = 32'd3272;
			62265: outdata = 32'd3271;
			62266: outdata = 32'd3270;
			62267: outdata = 32'd3269;
			62268: outdata = 32'd3268;
			62269: outdata = 32'd3267;
			62270: outdata = 32'd3266;
			62271: outdata = 32'd3265;
			62272: outdata = 32'd3264;
			62273: outdata = 32'd3263;
			62274: outdata = 32'd3262;
			62275: outdata = 32'd3261;
			62276: outdata = 32'd3260;
			62277: outdata = 32'd3259;
			62278: outdata = 32'd3258;
			62279: outdata = 32'd3257;
			62280: outdata = 32'd3256;
			62281: outdata = 32'd3255;
			62282: outdata = 32'd3254;
			62283: outdata = 32'd3253;
			62284: outdata = 32'd3252;
			62285: outdata = 32'd3251;
			62286: outdata = 32'd3250;
			62287: outdata = 32'd3249;
			62288: outdata = 32'd3248;
			62289: outdata = 32'd3247;
			62290: outdata = 32'd3246;
			62291: outdata = 32'd3245;
			62292: outdata = 32'd3244;
			62293: outdata = 32'd3243;
			62294: outdata = 32'd3242;
			62295: outdata = 32'd3241;
			62296: outdata = 32'd3240;
			62297: outdata = 32'd3239;
			62298: outdata = 32'd3238;
			62299: outdata = 32'd3237;
			62300: outdata = 32'd3236;
			62301: outdata = 32'd3235;
			62302: outdata = 32'd3234;
			62303: outdata = 32'd3233;
			62304: outdata = 32'd3232;
			62305: outdata = 32'd3231;
			62306: outdata = 32'd3230;
			62307: outdata = 32'd3229;
			62308: outdata = 32'd3228;
			62309: outdata = 32'd3227;
			62310: outdata = 32'd3226;
			62311: outdata = 32'd3225;
			62312: outdata = 32'd3224;
			62313: outdata = 32'd3223;
			62314: outdata = 32'd3222;
			62315: outdata = 32'd3221;
			62316: outdata = 32'd3220;
			62317: outdata = 32'd3219;
			62318: outdata = 32'd3218;
			62319: outdata = 32'd3217;
			62320: outdata = 32'd3216;
			62321: outdata = 32'd3215;
			62322: outdata = 32'd3214;
			62323: outdata = 32'd3213;
			62324: outdata = 32'd3212;
			62325: outdata = 32'd3211;
			62326: outdata = 32'd3210;
			62327: outdata = 32'd3209;
			62328: outdata = 32'd3208;
			62329: outdata = 32'd3207;
			62330: outdata = 32'd3206;
			62331: outdata = 32'd3205;
			62332: outdata = 32'd3204;
			62333: outdata = 32'd3203;
			62334: outdata = 32'd3202;
			62335: outdata = 32'd3201;
			62336: outdata = 32'd3200;
			62337: outdata = 32'd3199;
			62338: outdata = 32'd3198;
			62339: outdata = 32'd3197;
			62340: outdata = 32'd3196;
			62341: outdata = 32'd3195;
			62342: outdata = 32'd3194;
			62343: outdata = 32'd3193;
			62344: outdata = 32'd3192;
			62345: outdata = 32'd3191;
			62346: outdata = 32'd3190;
			62347: outdata = 32'd3189;
			62348: outdata = 32'd3188;
			62349: outdata = 32'd3187;
			62350: outdata = 32'd3186;
			62351: outdata = 32'd3185;
			62352: outdata = 32'd3184;
			62353: outdata = 32'd3183;
			62354: outdata = 32'd3182;
			62355: outdata = 32'd3181;
			62356: outdata = 32'd3180;
			62357: outdata = 32'd3179;
			62358: outdata = 32'd3178;
			62359: outdata = 32'd3177;
			62360: outdata = 32'd3176;
			62361: outdata = 32'd3175;
			62362: outdata = 32'd3174;
			62363: outdata = 32'd3173;
			62364: outdata = 32'd3172;
			62365: outdata = 32'd3171;
			62366: outdata = 32'd3170;
			62367: outdata = 32'd3169;
			62368: outdata = 32'd3168;
			62369: outdata = 32'd3167;
			62370: outdata = 32'd3166;
			62371: outdata = 32'd3165;
			62372: outdata = 32'd3164;
			62373: outdata = 32'd3163;
			62374: outdata = 32'd3162;
			62375: outdata = 32'd3161;
			62376: outdata = 32'd3160;
			62377: outdata = 32'd3159;
			62378: outdata = 32'd3158;
			62379: outdata = 32'd3157;
			62380: outdata = 32'd3156;
			62381: outdata = 32'd3155;
			62382: outdata = 32'd3154;
			62383: outdata = 32'd3153;
			62384: outdata = 32'd3152;
			62385: outdata = 32'd3151;
			62386: outdata = 32'd3150;
			62387: outdata = 32'd3149;
			62388: outdata = 32'd3148;
			62389: outdata = 32'd3147;
			62390: outdata = 32'd3146;
			62391: outdata = 32'd3145;
			62392: outdata = 32'd3144;
			62393: outdata = 32'd3143;
			62394: outdata = 32'd3142;
			62395: outdata = 32'd3141;
			62396: outdata = 32'd3140;
			62397: outdata = 32'd3139;
			62398: outdata = 32'd3138;
			62399: outdata = 32'd3137;
			62400: outdata = 32'd3136;
			62401: outdata = 32'd3135;
			62402: outdata = 32'd3134;
			62403: outdata = 32'd3133;
			62404: outdata = 32'd3132;
			62405: outdata = 32'd3131;
			62406: outdata = 32'd3130;
			62407: outdata = 32'd3129;
			62408: outdata = 32'd3128;
			62409: outdata = 32'd3127;
			62410: outdata = 32'd3126;
			62411: outdata = 32'd3125;
			62412: outdata = 32'd3124;
			62413: outdata = 32'd3123;
			62414: outdata = 32'd3122;
			62415: outdata = 32'd3121;
			62416: outdata = 32'd3120;
			62417: outdata = 32'd3119;
			62418: outdata = 32'd3118;
			62419: outdata = 32'd3117;
			62420: outdata = 32'd3116;
			62421: outdata = 32'd3115;
			62422: outdata = 32'd3114;
			62423: outdata = 32'd3113;
			62424: outdata = 32'd3112;
			62425: outdata = 32'd3111;
			62426: outdata = 32'd3110;
			62427: outdata = 32'd3109;
			62428: outdata = 32'd3108;
			62429: outdata = 32'd3107;
			62430: outdata = 32'd3106;
			62431: outdata = 32'd3105;
			62432: outdata = 32'd3104;
			62433: outdata = 32'd3103;
			62434: outdata = 32'd3102;
			62435: outdata = 32'd3101;
			62436: outdata = 32'd3100;
			62437: outdata = 32'd3099;
			62438: outdata = 32'd3098;
			62439: outdata = 32'd3097;
			62440: outdata = 32'd3096;
			62441: outdata = 32'd3095;
			62442: outdata = 32'd3094;
			62443: outdata = 32'd3093;
			62444: outdata = 32'd3092;
			62445: outdata = 32'd3091;
			62446: outdata = 32'd3090;
			62447: outdata = 32'd3089;
			62448: outdata = 32'd3088;
			62449: outdata = 32'd3087;
			62450: outdata = 32'd3086;
			62451: outdata = 32'd3085;
			62452: outdata = 32'd3084;
			62453: outdata = 32'd3083;
			62454: outdata = 32'd3082;
			62455: outdata = 32'd3081;
			62456: outdata = 32'd3080;
			62457: outdata = 32'd3079;
			62458: outdata = 32'd3078;
			62459: outdata = 32'd3077;
			62460: outdata = 32'd3076;
			62461: outdata = 32'd3075;
			62462: outdata = 32'd3074;
			62463: outdata = 32'd3073;
			62464: outdata = 32'd3072;
			62465: outdata = 32'd3071;
			62466: outdata = 32'd3070;
			62467: outdata = 32'd3069;
			62468: outdata = 32'd3068;
			62469: outdata = 32'd3067;
			62470: outdata = 32'd3066;
			62471: outdata = 32'd3065;
			62472: outdata = 32'd3064;
			62473: outdata = 32'd3063;
			62474: outdata = 32'd3062;
			62475: outdata = 32'd3061;
			62476: outdata = 32'd3060;
			62477: outdata = 32'd3059;
			62478: outdata = 32'd3058;
			62479: outdata = 32'd3057;
			62480: outdata = 32'd3056;
			62481: outdata = 32'd3055;
			62482: outdata = 32'd3054;
			62483: outdata = 32'd3053;
			62484: outdata = 32'd3052;
			62485: outdata = 32'd3051;
			62486: outdata = 32'd3050;
			62487: outdata = 32'd3049;
			62488: outdata = 32'd3048;
			62489: outdata = 32'd3047;
			62490: outdata = 32'd3046;
			62491: outdata = 32'd3045;
			62492: outdata = 32'd3044;
			62493: outdata = 32'd3043;
			62494: outdata = 32'd3042;
			62495: outdata = 32'd3041;
			62496: outdata = 32'd3040;
			62497: outdata = 32'd3039;
			62498: outdata = 32'd3038;
			62499: outdata = 32'd3037;
			62500: outdata = 32'd3036;
			62501: outdata = 32'd3035;
			62502: outdata = 32'd3034;
			62503: outdata = 32'd3033;
			62504: outdata = 32'd3032;
			62505: outdata = 32'd3031;
			62506: outdata = 32'd3030;
			62507: outdata = 32'd3029;
			62508: outdata = 32'd3028;
			62509: outdata = 32'd3027;
			62510: outdata = 32'd3026;
			62511: outdata = 32'd3025;
			62512: outdata = 32'd3024;
			62513: outdata = 32'd3023;
			62514: outdata = 32'd3022;
			62515: outdata = 32'd3021;
			62516: outdata = 32'd3020;
			62517: outdata = 32'd3019;
			62518: outdata = 32'd3018;
			62519: outdata = 32'd3017;
			62520: outdata = 32'd3016;
			62521: outdata = 32'd3015;
			62522: outdata = 32'd3014;
			62523: outdata = 32'd3013;
			62524: outdata = 32'd3012;
			62525: outdata = 32'd3011;
			62526: outdata = 32'd3010;
			62527: outdata = 32'd3009;
			62528: outdata = 32'd3008;
			62529: outdata = 32'd3007;
			62530: outdata = 32'd3006;
			62531: outdata = 32'd3005;
			62532: outdata = 32'd3004;
			62533: outdata = 32'd3003;
			62534: outdata = 32'd3002;
			62535: outdata = 32'd3001;
			62536: outdata = 32'd3000;
			62537: outdata = 32'd2999;
			62538: outdata = 32'd2998;
			62539: outdata = 32'd2997;
			62540: outdata = 32'd2996;
			62541: outdata = 32'd2995;
			62542: outdata = 32'd2994;
			62543: outdata = 32'd2993;
			62544: outdata = 32'd2992;
			62545: outdata = 32'd2991;
			62546: outdata = 32'd2990;
			62547: outdata = 32'd2989;
			62548: outdata = 32'd2988;
			62549: outdata = 32'd2987;
			62550: outdata = 32'd2986;
			62551: outdata = 32'd2985;
			62552: outdata = 32'd2984;
			62553: outdata = 32'd2983;
			62554: outdata = 32'd2982;
			62555: outdata = 32'd2981;
			62556: outdata = 32'd2980;
			62557: outdata = 32'd2979;
			62558: outdata = 32'd2978;
			62559: outdata = 32'd2977;
			62560: outdata = 32'd2976;
			62561: outdata = 32'd2975;
			62562: outdata = 32'd2974;
			62563: outdata = 32'd2973;
			62564: outdata = 32'd2972;
			62565: outdata = 32'd2971;
			62566: outdata = 32'd2970;
			62567: outdata = 32'd2969;
			62568: outdata = 32'd2968;
			62569: outdata = 32'd2967;
			62570: outdata = 32'd2966;
			62571: outdata = 32'd2965;
			62572: outdata = 32'd2964;
			62573: outdata = 32'd2963;
			62574: outdata = 32'd2962;
			62575: outdata = 32'd2961;
			62576: outdata = 32'd2960;
			62577: outdata = 32'd2959;
			62578: outdata = 32'd2958;
			62579: outdata = 32'd2957;
			62580: outdata = 32'd2956;
			62581: outdata = 32'd2955;
			62582: outdata = 32'd2954;
			62583: outdata = 32'd2953;
			62584: outdata = 32'd2952;
			62585: outdata = 32'd2951;
			62586: outdata = 32'd2950;
			62587: outdata = 32'd2949;
			62588: outdata = 32'd2948;
			62589: outdata = 32'd2947;
			62590: outdata = 32'd2946;
			62591: outdata = 32'd2945;
			62592: outdata = 32'd2944;
			62593: outdata = 32'd2943;
			62594: outdata = 32'd2942;
			62595: outdata = 32'd2941;
			62596: outdata = 32'd2940;
			62597: outdata = 32'd2939;
			62598: outdata = 32'd2938;
			62599: outdata = 32'd2937;
			62600: outdata = 32'd2936;
			62601: outdata = 32'd2935;
			62602: outdata = 32'd2934;
			62603: outdata = 32'd2933;
			62604: outdata = 32'd2932;
			62605: outdata = 32'd2931;
			62606: outdata = 32'd2930;
			62607: outdata = 32'd2929;
			62608: outdata = 32'd2928;
			62609: outdata = 32'd2927;
			62610: outdata = 32'd2926;
			62611: outdata = 32'd2925;
			62612: outdata = 32'd2924;
			62613: outdata = 32'd2923;
			62614: outdata = 32'd2922;
			62615: outdata = 32'd2921;
			62616: outdata = 32'd2920;
			62617: outdata = 32'd2919;
			62618: outdata = 32'd2918;
			62619: outdata = 32'd2917;
			62620: outdata = 32'd2916;
			62621: outdata = 32'd2915;
			62622: outdata = 32'd2914;
			62623: outdata = 32'd2913;
			62624: outdata = 32'd2912;
			62625: outdata = 32'd2911;
			62626: outdata = 32'd2910;
			62627: outdata = 32'd2909;
			62628: outdata = 32'd2908;
			62629: outdata = 32'd2907;
			62630: outdata = 32'd2906;
			62631: outdata = 32'd2905;
			62632: outdata = 32'd2904;
			62633: outdata = 32'd2903;
			62634: outdata = 32'd2902;
			62635: outdata = 32'd2901;
			62636: outdata = 32'd2900;
			62637: outdata = 32'd2899;
			62638: outdata = 32'd2898;
			62639: outdata = 32'd2897;
			62640: outdata = 32'd2896;
			62641: outdata = 32'd2895;
			62642: outdata = 32'd2894;
			62643: outdata = 32'd2893;
			62644: outdata = 32'd2892;
			62645: outdata = 32'd2891;
			62646: outdata = 32'd2890;
			62647: outdata = 32'd2889;
			62648: outdata = 32'd2888;
			62649: outdata = 32'd2887;
			62650: outdata = 32'd2886;
			62651: outdata = 32'd2885;
			62652: outdata = 32'd2884;
			62653: outdata = 32'd2883;
			62654: outdata = 32'd2882;
			62655: outdata = 32'd2881;
			62656: outdata = 32'd2880;
			62657: outdata = 32'd2879;
			62658: outdata = 32'd2878;
			62659: outdata = 32'd2877;
			62660: outdata = 32'd2876;
			62661: outdata = 32'd2875;
			62662: outdata = 32'd2874;
			62663: outdata = 32'd2873;
			62664: outdata = 32'd2872;
			62665: outdata = 32'd2871;
			62666: outdata = 32'd2870;
			62667: outdata = 32'd2869;
			62668: outdata = 32'd2868;
			62669: outdata = 32'd2867;
			62670: outdata = 32'd2866;
			62671: outdata = 32'd2865;
			62672: outdata = 32'd2864;
			62673: outdata = 32'd2863;
			62674: outdata = 32'd2862;
			62675: outdata = 32'd2861;
			62676: outdata = 32'd2860;
			62677: outdata = 32'd2859;
			62678: outdata = 32'd2858;
			62679: outdata = 32'd2857;
			62680: outdata = 32'd2856;
			62681: outdata = 32'd2855;
			62682: outdata = 32'd2854;
			62683: outdata = 32'd2853;
			62684: outdata = 32'd2852;
			62685: outdata = 32'd2851;
			62686: outdata = 32'd2850;
			62687: outdata = 32'd2849;
			62688: outdata = 32'd2848;
			62689: outdata = 32'd2847;
			62690: outdata = 32'd2846;
			62691: outdata = 32'd2845;
			62692: outdata = 32'd2844;
			62693: outdata = 32'd2843;
			62694: outdata = 32'd2842;
			62695: outdata = 32'd2841;
			62696: outdata = 32'd2840;
			62697: outdata = 32'd2839;
			62698: outdata = 32'd2838;
			62699: outdata = 32'd2837;
			62700: outdata = 32'd2836;
			62701: outdata = 32'd2835;
			62702: outdata = 32'd2834;
			62703: outdata = 32'd2833;
			62704: outdata = 32'd2832;
			62705: outdata = 32'd2831;
			62706: outdata = 32'd2830;
			62707: outdata = 32'd2829;
			62708: outdata = 32'd2828;
			62709: outdata = 32'd2827;
			62710: outdata = 32'd2826;
			62711: outdata = 32'd2825;
			62712: outdata = 32'd2824;
			62713: outdata = 32'd2823;
			62714: outdata = 32'd2822;
			62715: outdata = 32'd2821;
			62716: outdata = 32'd2820;
			62717: outdata = 32'd2819;
			62718: outdata = 32'd2818;
			62719: outdata = 32'd2817;
			62720: outdata = 32'd2816;
			62721: outdata = 32'd2815;
			62722: outdata = 32'd2814;
			62723: outdata = 32'd2813;
			62724: outdata = 32'd2812;
			62725: outdata = 32'd2811;
			62726: outdata = 32'd2810;
			62727: outdata = 32'd2809;
			62728: outdata = 32'd2808;
			62729: outdata = 32'd2807;
			62730: outdata = 32'd2806;
			62731: outdata = 32'd2805;
			62732: outdata = 32'd2804;
			62733: outdata = 32'd2803;
			62734: outdata = 32'd2802;
			62735: outdata = 32'd2801;
			62736: outdata = 32'd2800;
			62737: outdata = 32'd2799;
			62738: outdata = 32'd2798;
			62739: outdata = 32'd2797;
			62740: outdata = 32'd2796;
			62741: outdata = 32'd2795;
			62742: outdata = 32'd2794;
			62743: outdata = 32'd2793;
			62744: outdata = 32'd2792;
			62745: outdata = 32'd2791;
			62746: outdata = 32'd2790;
			62747: outdata = 32'd2789;
			62748: outdata = 32'd2788;
			62749: outdata = 32'd2787;
			62750: outdata = 32'd2786;
			62751: outdata = 32'd2785;
			62752: outdata = 32'd2784;
			62753: outdata = 32'd2783;
			62754: outdata = 32'd2782;
			62755: outdata = 32'd2781;
			62756: outdata = 32'd2780;
			62757: outdata = 32'd2779;
			62758: outdata = 32'd2778;
			62759: outdata = 32'd2777;
			62760: outdata = 32'd2776;
			62761: outdata = 32'd2775;
			62762: outdata = 32'd2774;
			62763: outdata = 32'd2773;
			62764: outdata = 32'd2772;
			62765: outdata = 32'd2771;
			62766: outdata = 32'd2770;
			62767: outdata = 32'd2769;
			62768: outdata = 32'd2768;
			62769: outdata = 32'd2767;
			62770: outdata = 32'd2766;
			62771: outdata = 32'd2765;
			62772: outdata = 32'd2764;
			62773: outdata = 32'd2763;
			62774: outdata = 32'd2762;
			62775: outdata = 32'd2761;
			62776: outdata = 32'd2760;
			62777: outdata = 32'd2759;
			62778: outdata = 32'd2758;
			62779: outdata = 32'd2757;
			62780: outdata = 32'd2756;
			62781: outdata = 32'd2755;
			62782: outdata = 32'd2754;
			62783: outdata = 32'd2753;
			62784: outdata = 32'd2752;
			62785: outdata = 32'd2751;
			62786: outdata = 32'd2750;
			62787: outdata = 32'd2749;
			62788: outdata = 32'd2748;
			62789: outdata = 32'd2747;
			62790: outdata = 32'd2746;
			62791: outdata = 32'd2745;
			62792: outdata = 32'd2744;
			62793: outdata = 32'd2743;
			62794: outdata = 32'd2742;
			62795: outdata = 32'd2741;
			62796: outdata = 32'd2740;
			62797: outdata = 32'd2739;
			62798: outdata = 32'd2738;
			62799: outdata = 32'd2737;
			62800: outdata = 32'd2736;
			62801: outdata = 32'd2735;
			62802: outdata = 32'd2734;
			62803: outdata = 32'd2733;
			62804: outdata = 32'd2732;
			62805: outdata = 32'd2731;
			62806: outdata = 32'd2730;
			62807: outdata = 32'd2729;
			62808: outdata = 32'd2728;
			62809: outdata = 32'd2727;
			62810: outdata = 32'd2726;
			62811: outdata = 32'd2725;
			62812: outdata = 32'd2724;
			62813: outdata = 32'd2723;
			62814: outdata = 32'd2722;
			62815: outdata = 32'd2721;
			62816: outdata = 32'd2720;
			62817: outdata = 32'd2719;
			62818: outdata = 32'd2718;
			62819: outdata = 32'd2717;
			62820: outdata = 32'd2716;
			62821: outdata = 32'd2715;
			62822: outdata = 32'd2714;
			62823: outdata = 32'd2713;
			62824: outdata = 32'd2712;
			62825: outdata = 32'd2711;
			62826: outdata = 32'd2710;
			62827: outdata = 32'd2709;
			62828: outdata = 32'd2708;
			62829: outdata = 32'd2707;
			62830: outdata = 32'd2706;
			62831: outdata = 32'd2705;
			62832: outdata = 32'd2704;
			62833: outdata = 32'd2703;
			62834: outdata = 32'd2702;
			62835: outdata = 32'd2701;
			62836: outdata = 32'd2700;
			62837: outdata = 32'd2699;
			62838: outdata = 32'd2698;
			62839: outdata = 32'd2697;
			62840: outdata = 32'd2696;
			62841: outdata = 32'd2695;
			62842: outdata = 32'd2694;
			62843: outdata = 32'd2693;
			62844: outdata = 32'd2692;
			62845: outdata = 32'd2691;
			62846: outdata = 32'd2690;
			62847: outdata = 32'd2689;
			62848: outdata = 32'd2688;
			62849: outdata = 32'd2687;
			62850: outdata = 32'd2686;
			62851: outdata = 32'd2685;
			62852: outdata = 32'd2684;
			62853: outdata = 32'd2683;
			62854: outdata = 32'd2682;
			62855: outdata = 32'd2681;
			62856: outdata = 32'd2680;
			62857: outdata = 32'd2679;
			62858: outdata = 32'd2678;
			62859: outdata = 32'd2677;
			62860: outdata = 32'd2676;
			62861: outdata = 32'd2675;
			62862: outdata = 32'd2674;
			62863: outdata = 32'd2673;
			62864: outdata = 32'd2672;
			62865: outdata = 32'd2671;
			62866: outdata = 32'd2670;
			62867: outdata = 32'd2669;
			62868: outdata = 32'd2668;
			62869: outdata = 32'd2667;
			62870: outdata = 32'd2666;
			62871: outdata = 32'd2665;
			62872: outdata = 32'd2664;
			62873: outdata = 32'd2663;
			62874: outdata = 32'd2662;
			62875: outdata = 32'd2661;
			62876: outdata = 32'd2660;
			62877: outdata = 32'd2659;
			62878: outdata = 32'd2658;
			62879: outdata = 32'd2657;
			62880: outdata = 32'd2656;
			62881: outdata = 32'd2655;
			62882: outdata = 32'd2654;
			62883: outdata = 32'd2653;
			62884: outdata = 32'd2652;
			62885: outdata = 32'd2651;
			62886: outdata = 32'd2650;
			62887: outdata = 32'd2649;
			62888: outdata = 32'd2648;
			62889: outdata = 32'd2647;
			62890: outdata = 32'd2646;
			62891: outdata = 32'd2645;
			62892: outdata = 32'd2644;
			62893: outdata = 32'd2643;
			62894: outdata = 32'd2642;
			62895: outdata = 32'd2641;
			62896: outdata = 32'd2640;
			62897: outdata = 32'd2639;
			62898: outdata = 32'd2638;
			62899: outdata = 32'd2637;
			62900: outdata = 32'd2636;
			62901: outdata = 32'd2635;
			62902: outdata = 32'd2634;
			62903: outdata = 32'd2633;
			62904: outdata = 32'd2632;
			62905: outdata = 32'd2631;
			62906: outdata = 32'd2630;
			62907: outdata = 32'd2629;
			62908: outdata = 32'd2628;
			62909: outdata = 32'd2627;
			62910: outdata = 32'd2626;
			62911: outdata = 32'd2625;
			62912: outdata = 32'd2624;
			62913: outdata = 32'd2623;
			62914: outdata = 32'd2622;
			62915: outdata = 32'd2621;
			62916: outdata = 32'd2620;
			62917: outdata = 32'd2619;
			62918: outdata = 32'd2618;
			62919: outdata = 32'd2617;
			62920: outdata = 32'd2616;
			62921: outdata = 32'd2615;
			62922: outdata = 32'd2614;
			62923: outdata = 32'd2613;
			62924: outdata = 32'd2612;
			62925: outdata = 32'd2611;
			62926: outdata = 32'd2610;
			62927: outdata = 32'd2609;
			62928: outdata = 32'd2608;
			62929: outdata = 32'd2607;
			62930: outdata = 32'd2606;
			62931: outdata = 32'd2605;
			62932: outdata = 32'd2604;
			62933: outdata = 32'd2603;
			62934: outdata = 32'd2602;
			62935: outdata = 32'd2601;
			62936: outdata = 32'd2600;
			62937: outdata = 32'd2599;
			62938: outdata = 32'd2598;
			62939: outdata = 32'd2597;
			62940: outdata = 32'd2596;
			62941: outdata = 32'd2595;
			62942: outdata = 32'd2594;
			62943: outdata = 32'd2593;
			62944: outdata = 32'd2592;
			62945: outdata = 32'd2591;
			62946: outdata = 32'd2590;
			62947: outdata = 32'd2589;
			62948: outdata = 32'd2588;
			62949: outdata = 32'd2587;
			62950: outdata = 32'd2586;
			62951: outdata = 32'd2585;
			62952: outdata = 32'd2584;
			62953: outdata = 32'd2583;
			62954: outdata = 32'd2582;
			62955: outdata = 32'd2581;
			62956: outdata = 32'd2580;
			62957: outdata = 32'd2579;
			62958: outdata = 32'd2578;
			62959: outdata = 32'd2577;
			62960: outdata = 32'd2576;
			62961: outdata = 32'd2575;
			62962: outdata = 32'd2574;
			62963: outdata = 32'd2573;
			62964: outdata = 32'd2572;
			62965: outdata = 32'd2571;
			62966: outdata = 32'd2570;
			62967: outdata = 32'd2569;
			62968: outdata = 32'd2568;
			62969: outdata = 32'd2567;
			62970: outdata = 32'd2566;
			62971: outdata = 32'd2565;
			62972: outdata = 32'd2564;
			62973: outdata = 32'd2563;
			62974: outdata = 32'd2562;
			62975: outdata = 32'd2561;
			62976: outdata = 32'd2560;
			62977: outdata = 32'd2559;
			62978: outdata = 32'd2558;
			62979: outdata = 32'd2557;
			62980: outdata = 32'd2556;
			62981: outdata = 32'd2555;
			62982: outdata = 32'd2554;
			62983: outdata = 32'd2553;
			62984: outdata = 32'd2552;
			62985: outdata = 32'd2551;
			62986: outdata = 32'd2550;
			62987: outdata = 32'd2549;
			62988: outdata = 32'd2548;
			62989: outdata = 32'd2547;
			62990: outdata = 32'd2546;
			62991: outdata = 32'd2545;
			62992: outdata = 32'd2544;
			62993: outdata = 32'd2543;
			62994: outdata = 32'd2542;
			62995: outdata = 32'd2541;
			62996: outdata = 32'd2540;
			62997: outdata = 32'd2539;
			62998: outdata = 32'd2538;
			62999: outdata = 32'd2537;
			63000: outdata = 32'd2536;
			63001: outdata = 32'd2535;
			63002: outdata = 32'd2534;
			63003: outdata = 32'd2533;
			63004: outdata = 32'd2532;
			63005: outdata = 32'd2531;
			63006: outdata = 32'd2530;
			63007: outdata = 32'd2529;
			63008: outdata = 32'd2528;
			63009: outdata = 32'd2527;
			63010: outdata = 32'd2526;
			63011: outdata = 32'd2525;
			63012: outdata = 32'd2524;
			63013: outdata = 32'd2523;
			63014: outdata = 32'd2522;
			63015: outdata = 32'd2521;
			63016: outdata = 32'd2520;
			63017: outdata = 32'd2519;
			63018: outdata = 32'd2518;
			63019: outdata = 32'd2517;
			63020: outdata = 32'd2516;
			63021: outdata = 32'd2515;
			63022: outdata = 32'd2514;
			63023: outdata = 32'd2513;
			63024: outdata = 32'd2512;
			63025: outdata = 32'd2511;
			63026: outdata = 32'd2510;
			63027: outdata = 32'd2509;
			63028: outdata = 32'd2508;
			63029: outdata = 32'd2507;
			63030: outdata = 32'd2506;
			63031: outdata = 32'd2505;
			63032: outdata = 32'd2504;
			63033: outdata = 32'd2503;
			63034: outdata = 32'd2502;
			63035: outdata = 32'd2501;
			63036: outdata = 32'd2500;
			63037: outdata = 32'd2499;
			63038: outdata = 32'd2498;
			63039: outdata = 32'd2497;
			63040: outdata = 32'd2496;
			63041: outdata = 32'd2495;
			63042: outdata = 32'd2494;
			63043: outdata = 32'd2493;
			63044: outdata = 32'd2492;
			63045: outdata = 32'd2491;
			63046: outdata = 32'd2490;
			63047: outdata = 32'd2489;
			63048: outdata = 32'd2488;
			63049: outdata = 32'd2487;
			63050: outdata = 32'd2486;
			63051: outdata = 32'd2485;
			63052: outdata = 32'd2484;
			63053: outdata = 32'd2483;
			63054: outdata = 32'd2482;
			63055: outdata = 32'd2481;
			63056: outdata = 32'd2480;
			63057: outdata = 32'd2479;
			63058: outdata = 32'd2478;
			63059: outdata = 32'd2477;
			63060: outdata = 32'd2476;
			63061: outdata = 32'd2475;
			63062: outdata = 32'd2474;
			63063: outdata = 32'd2473;
			63064: outdata = 32'd2472;
			63065: outdata = 32'd2471;
			63066: outdata = 32'd2470;
			63067: outdata = 32'd2469;
			63068: outdata = 32'd2468;
			63069: outdata = 32'd2467;
			63070: outdata = 32'd2466;
			63071: outdata = 32'd2465;
			63072: outdata = 32'd2464;
			63073: outdata = 32'd2463;
			63074: outdata = 32'd2462;
			63075: outdata = 32'd2461;
			63076: outdata = 32'd2460;
			63077: outdata = 32'd2459;
			63078: outdata = 32'd2458;
			63079: outdata = 32'd2457;
			63080: outdata = 32'd2456;
			63081: outdata = 32'd2455;
			63082: outdata = 32'd2454;
			63083: outdata = 32'd2453;
			63084: outdata = 32'd2452;
			63085: outdata = 32'd2451;
			63086: outdata = 32'd2450;
			63087: outdata = 32'd2449;
			63088: outdata = 32'd2448;
			63089: outdata = 32'd2447;
			63090: outdata = 32'd2446;
			63091: outdata = 32'd2445;
			63092: outdata = 32'd2444;
			63093: outdata = 32'd2443;
			63094: outdata = 32'd2442;
			63095: outdata = 32'd2441;
			63096: outdata = 32'd2440;
			63097: outdata = 32'd2439;
			63098: outdata = 32'd2438;
			63099: outdata = 32'd2437;
			63100: outdata = 32'd2436;
			63101: outdata = 32'd2435;
			63102: outdata = 32'd2434;
			63103: outdata = 32'd2433;
			63104: outdata = 32'd2432;
			63105: outdata = 32'd2431;
			63106: outdata = 32'd2430;
			63107: outdata = 32'd2429;
			63108: outdata = 32'd2428;
			63109: outdata = 32'd2427;
			63110: outdata = 32'd2426;
			63111: outdata = 32'd2425;
			63112: outdata = 32'd2424;
			63113: outdata = 32'd2423;
			63114: outdata = 32'd2422;
			63115: outdata = 32'd2421;
			63116: outdata = 32'd2420;
			63117: outdata = 32'd2419;
			63118: outdata = 32'd2418;
			63119: outdata = 32'd2417;
			63120: outdata = 32'd2416;
			63121: outdata = 32'd2415;
			63122: outdata = 32'd2414;
			63123: outdata = 32'd2413;
			63124: outdata = 32'd2412;
			63125: outdata = 32'd2411;
			63126: outdata = 32'd2410;
			63127: outdata = 32'd2409;
			63128: outdata = 32'd2408;
			63129: outdata = 32'd2407;
			63130: outdata = 32'd2406;
			63131: outdata = 32'd2405;
			63132: outdata = 32'd2404;
			63133: outdata = 32'd2403;
			63134: outdata = 32'd2402;
			63135: outdata = 32'd2401;
			63136: outdata = 32'd2400;
			63137: outdata = 32'd2399;
			63138: outdata = 32'd2398;
			63139: outdata = 32'd2397;
			63140: outdata = 32'd2396;
			63141: outdata = 32'd2395;
			63142: outdata = 32'd2394;
			63143: outdata = 32'd2393;
			63144: outdata = 32'd2392;
			63145: outdata = 32'd2391;
			63146: outdata = 32'd2390;
			63147: outdata = 32'd2389;
			63148: outdata = 32'd2388;
			63149: outdata = 32'd2387;
			63150: outdata = 32'd2386;
			63151: outdata = 32'd2385;
			63152: outdata = 32'd2384;
			63153: outdata = 32'd2383;
			63154: outdata = 32'd2382;
			63155: outdata = 32'd2381;
			63156: outdata = 32'd2380;
			63157: outdata = 32'd2379;
			63158: outdata = 32'd2378;
			63159: outdata = 32'd2377;
			63160: outdata = 32'd2376;
			63161: outdata = 32'd2375;
			63162: outdata = 32'd2374;
			63163: outdata = 32'd2373;
			63164: outdata = 32'd2372;
			63165: outdata = 32'd2371;
			63166: outdata = 32'd2370;
			63167: outdata = 32'd2369;
			63168: outdata = 32'd2368;
			63169: outdata = 32'd2367;
			63170: outdata = 32'd2366;
			63171: outdata = 32'd2365;
			63172: outdata = 32'd2364;
			63173: outdata = 32'd2363;
			63174: outdata = 32'd2362;
			63175: outdata = 32'd2361;
			63176: outdata = 32'd2360;
			63177: outdata = 32'd2359;
			63178: outdata = 32'd2358;
			63179: outdata = 32'd2357;
			63180: outdata = 32'd2356;
			63181: outdata = 32'd2355;
			63182: outdata = 32'd2354;
			63183: outdata = 32'd2353;
			63184: outdata = 32'd2352;
			63185: outdata = 32'd2351;
			63186: outdata = 32'd2350;
			63187: outdata = 32'd2349;
			63188: outdata = 32'd2348;
			63189: outdata = 32'd2347;
			63190: outdata = 32'd2346;
			63191: outdata = 32'd2345;
			63192: outdata = 32'd2344;
			63193: outdata = 32'd2343;
			63194: outdata = 32'd2342;
			63195: outdata = 32'd2341;
			63196: outdata = 32'd2340;
			63197: outdata = 32'd2339;
			63198: outdata = 32'd2338;
			63199: outdata = 32'd2337;
			63200: outdata = 32'd2336;
			63201: outdata = 32'd2335;
			63202: outdata = 32'd2334;
			63203: outdata = 32'd2333;
			63204: outdata = 32'd2332;
			63205: outdata = 32'd2331;
			63206: outdata = 32'd2330;
			63207: outdata = 32'd2329;
			63208: outdata = 32'd2328;
			63209: outdata = 32'd2327;
			63210: outdata = 32'd2326;
			63211: outdata = 32'd2325;
			63212: outdata = 32'd2324;
			63213: outdata = 32'd2323;
			63214: outdata = 32'd2322;
			63215: outdata = 32'd2321;
			63216: outdata = 32'd2320;
			63217: outdata = 32'd2319;
			63218: outdata = 32'd2318;
			63219: outdata = 32'd2317;
			63220: outdata = 32'd2316;
			63221: outdata = 32'd2315;
			63222: outdata = 32'd2314;
			63223: outdata = 32'd2313;
			63224: outdata = 32'd2312;
			63225: outdata = 32'd2311;
			63226: outdata = 32'd2310;
			63227: outdata = 32'd2309;
			63228: outdata = 32'd2308;
			63229: outdata = 32'd2307;
			63230: outdata = 32'd2306;
			63231: outdata = 32'd2305;
			63232: outdata = 32'd2304;
			63233: outdata = 32'd2303;
			63234: outdata = 32'd2302;
			63235: outdata = 32'd2301;
			63236: outdata = 32'd2300;
			63237: outdata = 32'd2299;
			63238: outdata = 32'd2298;
			63239: outdata = 32'd2297;
			63240: outdata = 32'd2296;
			63241: outdata = 32'd2295;
			63242: outdata = 32'd2294;
			63243: outdata = 32'd2293;
			63244: outdata = 32'd2292;
			63245: outdata = 32'd2291;
			63246: outdata = 32'd2290;
			63247: outdata = 32'd2289;
			63248: outdata = 32'd2288;
			63249: outdata = 32'd2287;
			63250: outdata = 32'd2286;
			63251: outdata = 32'd2285;
			63252: outdata = 32'd2284;
			63253: outdata = 32'd2283;
			63254: outdata = 32'd2282;
			63255: outdata = 32'd2281;
			63256: outdata = 32'd2280;
			63257: outdata = 32'd2279;
			63258: outdata = 32'd2278;
			63259: outdata = 32'd2277;
			63260: outdata = 32'd2276;
			63261: outdata = 32'd2275;
			63262: outdata = 32'd2274;
			63263: outdata = 32'd2273;
			63264: outdata = 32'd2272;
			63265: outdata = 32'd2271;
			63266: outdata = 32'd2270;
			63267: outdata = 32'd2269;
			63268: outdata = 32'd2268;
			63269: outdata = 32'd2267;
			63270: outdata = 32'd2266;
			63271: outdata = 32'd2265;
			63272: outdata = 32'd2264;
			63273: outdata = 32'd2263;
			63274: outdata = 32'd2262;
			63275: outdata = 32'd2261;
			63276: outdata = 32'd2260;
			63277: outdata = 32'd2259;
			63278: outdata = 32'd2258;
			63279: outdata = 32'd2257;
			63280: outdata = 32'd2256;
			63281: outdata = 32'd2255;
			63282: outdata = 32'd2254;
			63283: outdata = 32'd2253;
			63284: outdata = 32'd2252;
			63285: outdata = 32'd2251;
			63286: outdata = 32'd2250;
			63287: outdata = 32'd2249;
			63288: outdata = 32'd2248;
			63289: outdata = 32'd2247;
			63290: outdata = 32'd2246;
			63291: outdata = 32'd2245;
			63292: outdata = 32'd2244;
			63293: outdata = 32'd2243;
			63294: outdata = 32'd2242;
			63295: outdata = 32'd2241;
			63296: outdata = 32'd2240;
			63297: outdata = 32'd2239;
			63298: outdata = 32'd2238;
			63299: outdata = 32'd2237;
			63300: outdata = 32'd2236;
			63301: outdata = 32'd2235;
			63302: outdata = 32'd2234;
			63303: outdata = 32'd2233;
			63304: outdata = 32'd2232;
			63305: outdata = 32'd2231;
			63306: outdata = 32'd2230;
			63307: outdata = 32'd2229;
			63308: outdata = 32'd2228;
			63309: outdata = 32'd2227;
			63310: outdata = 32'd2226;
			63311: outdata = 32'd2225;
			63312: outdata = 32'd2224;
			63313: outdata = 32'd2223;
			63314: outdata = 32'd2222;
			63315: outdata = 32'd2221;
			63316: outdata = 32'd2220;
			63317: outdata = 32'd2219;
			63318: outdata = 32'd2218;
			63319: outdata = 32'd2217;
			63320: outdata = 32'd2216;
			63321: outdata = 32'd2215;
			63322: outdata = 32'd2214;
			63323: outdata = 32'd2213;
			63324: outdata = 32'd2212;
			63325: outdata = 32'd2211;
			63326: outdata = 32'd2210;
			63327: outdata = 32'd2209;
			63328: outdata = 32'd2208;
			63329: outdata = 32'd2207;
			63330: outdata = 32'd2206;
			63331: outdata = 32'd2205;
			63332: outdata = 32'd2204;
			63333: outdata = 32'd2203;
			63334: outdata = 32'd2202;
			63335: outdata = 32'd2201;
			63336: outdata = 32'd2200;
			63337: outdata = 32'd2199;
			63338: outdata = 32'd2198;
			63339: outdata = 32'd2197;
			63340: outdata = 32'd2196;
			63341: outdata = 32'd2195;
			63342: outdata = 32'd2194;
			63343: outdata = 32'd2193;
			63344: outdata = 32'd2192;
			63345: outdata = 32'd2191;
			63346: outdata = 32'd2190;
			63347: outdata = 32'd2189;
			63348: outdata = 32'd2188;
			63349: outdata = 32'd2187;
			63350: outdata = 32'd2186;
			63351: outdata = 32'd2185;
			63352: outdata = 32'd2184;
			63353: outdata = 32'd2183;
			63354: outdata = 32'd2182;
			63355: outdata = 32'd2181;
			63356: outdata = 32'd2180;
			63357: outdata = 32'd2179;
			63358: outdata = 32'd2178;
			63359: outdata = 32'd2177;
			63360: outdata = 32'd2176;
			63361: outdata = 32'd2175;
			63362: outdata = 32'd2174;
			63363: outdata = 32'd2173;
			63364: outdata = 32'd2172;
			63365: outdata = 32'd2171;
			63366: outdata = 32'd2170;
			63367: outdata = 32'd2169;
			63368: outdata = 32'd2168;
			63369: outdata = 32'd2167;
			63370: outdata = 32'd2166;
			63371: outdata = 32'd2165;
			63372: outdata = 32'd2164;
			63373: outdata = 32'd2163;
			63374: outdata = 32'd2162;
			63375: outdata = 32'd2161;
			63376: outdata = 32'd2160;
			63377: outdata = 32'd2159;
			63378: outdata = 32'd2158;
			63379: outdata = 32'd2157;
			63380: outdata = 32'd2156;
			63381: outdata = 32'd2155;
			63382: outdata = 32'd2154;
			63383: outdata = 32'd2153;
			63384: outdata = 32'd2152;
			63385: outdata = 32'd2151;
			63386: outdata = 32'd2150;
			63387: outdata = 32'd2149;
			63388: outdata = 32'd2148;
			63389: outdata = 32'd2147;
			63390: outdata = 32'd2146;
			63391: outdata = 32'd2145;
			63392: outdata = 32'd2144;
			63393: outdata = 32'd2143;
			63394: outdata = 32'd2142;
			63395: outdata = 32'd2141;
			63396: outdata = 32'd2140;
			63397: outdata = 32'd2139;
			63398: outdata = 32'd2138;
			63399: outdata = 32'd2137;
			63400: outdata = 32'd2136;
			63401: outdata = 32'd2135;
			63402: outdata = 32'd2134;
			63403: outdata = 32'd2133;
			63404: outdata = 32'd2132;
			63405: outdata = 32'd2131;
			63406: outdata = 32'd2130;
			63407: outdata = 32'd2129;
			63408: outdata = 32'd2128;
			63409: outdata = 32'd2127;
			63410: outdata = 32'd2126;
			63411: outdata = 32'd2125;
			63412: outdata = 32'd2124;
			63413: outdata = 32'd2123;
			63414: outdata = 32'd2122;
			63415: outdata = 32'd2121;
			63416: outdata = 32'd2120;
			63417: outdata = 32'd2119;
			63418: outdata = 32'd2118;
			63419: outdata = 32'd2117;
			63420: outdata = 32'd2116;
			63421: outdata = 32'd2115;
			63422: outdata = 32'd2114;
			63423: outdata = 32'd2113;
			63424: outdata = 32'd2112;
			63425: outdata = 32'd2111;
			63426: outdata = 32'd2110;
			63427: outdata = 32'd2109;
			63428: outdata = 32'd2108;
			63429: outdata = 32'd2107;
			63430: outdata = 32'd2106;
			63431: outdata = 32'd2105;
			63432: outdata = 32'd2104;
			63433: outdata = 32'd2103;
			63434: outdata = 32'd2102;
			63435: outdata = 32'd2101;
			63436: outdata = 32'd2100;
			63437: outdata = 32'd2099;
			63438: outdata = 32'd2098;
			63439: outdata = 32'd2097;
			63440: outdata = 32'd2096;
			63441: outdata = 32'd2095;
			63442: outdata = 32'd2094;
			63443: outdata = 32'd2093;
			63444: outdata = 32'd2092;
			63445: outdata = 32'd2091;
			63446: outdata = 32'd2090;
			63447: outdata = 32'd2089;
			63448: outdata = 32'd2088;
			63449: outdata = 32'd2087;
			63450: outdata = 32'd2086;
			63451: outdata = 32'd2085;
			63452: outdata = 32'd2084;
			63453: outdata = 32'd2083;
			63454: outdata = 32'd2082;
			63455: outdata = 32'd2081;
			63456: outdata = 32'd2080;
			63457: outdata = 32'd2079;
			63458: outdata = 32'd2078;
			63459: outdata = 32'd2077;
			63460: outdata = 32'd2076;
			63461: outdata = 32'd2075;
			63462: outdata = 32'd2074;
			63463: outdata = 32'd2073;
			63464: outdata = 32'd2072;
			63465: outdata = 32'd2071;
			63466: outdata = 32'd2070;
			63467: outdata = 32'd2069;
			63468: outdata = 32'd2068;
			63469: outdata = 32'd2067;
			63470: outdata = 32'd2066;
			63471: outdata = 32'd2065;
			63472: outdata = 32'd2064;
			63473: outdata = 32'd2063;
			63474: outdata = 32'd2062;
			63475: outdata = 32'd2061;
			63476: outdata = 32'd2060;
			63477: outdata = 32'd2059;
			63478: outdata = 32'd2058;
			63479: outdata = 32'd2057;
			63480: outdata = 32'd2056;
			63481: outdata = 32'd2055;
			63482: outdata = 32'd2054;
			63483: outdata = 32'd2053;
			63484: outdata = 32'd2052;
			63485: outdata = 32'd2051;
			63486: outdata = 32'd2050;
			63487: outdata = 32'd2049;
			63488: outdata = 32'd2048;
			63489: outdata = 32'd2047;
			63490: outdata = 32'd2046;
			63491: outdata = 32'd2045;
			63492: outdata = 32'd2044;
			63493: outdata = 32'd2043;
			63494: outdata = 32'd2042;
			63495: outdata = 32'd2041;
			63496: outdata = 32'd2040;
			63497: outdata = 32'd2039;
			63498: outdata = 32'd2038;
			63499: outdata = 32'd2037;
			63500: outdata = 32'd2036;
			63501: outdata = 32'd2035;
			63502: outdata = 32'd2034;
			63503: outdata = 32'd2033;
			63504: outdata = 32'd2032;
			63505: outdata = 32'd2031;
			63506: outdata = 32'd2030;
			63507: outdata = 32'd2029;
			63508: outdata = 32'd2028;
			63509: outdata = 32'd2027;
			63510: outdata = 32'd2026;
			63511: outdata = 32'd2025;
			63512: outdata = 32'd2024;
			63513: outdata = 32'd2023;
			63514: outdata = 32'd2022;
			63515: outdata = 32'd2021;
			63516: outdata = 32'd2020;
			63517: outdata = 32'd2019;
			63518: outdata = 32'd2018;
			63519: outdata = 32'd2017;
			63520: outdata = 32'd2016;
			63521: outdata = 32'd2015;
			63522: outdata = 32'd2014;
			63523: outdata = 32'd2013;
			63524: outdata = 32'd2012;
			63525: outdata = 32'd2011;
			63526: outdata = 32'd2010;
			63527: outdata = 32'd2009;
			63528: outdata = 32'd2008;
			63529: outdata = 32'd2007;
			63530: outdata = 32'd2006;
			63531: outdata = 32'd2005;
			63532: outdata = 32'd2004;
			63533: outdata = 32'd2003;
			63534: outdata = 32'd2002;
			63535: outdata = 32'd2001;
			63536: outdata = 32'd2000;
			63537: outdata = 32'd1999;
			63538: outdata = 32'd1998;
			63539: outdata = 32'd1997;
			63540: outdata = 32'd1996;
			63541: outdata = 32'd1995;
			63542: outdata = 32'd1994;
			63543: outdata = 32'd1993;
			63544: outdata = 32'd1992;
			63545: outdata = 32'd1991;
			63546: outdata = 32'd1990;
			63547: outdata = 32'd1989;
			63548: outdata = 32'd1988;
			63549: outdata = 32'd1987;
			63550: outdata = 32'd1986;
			63551: outdata = 32'd1985;
			63552: outdata = 32'd1984;
			63553: outdata = 32'd1983;
			63554: outdata = 32'd1982;
			63555: outdata = 32'd1981;
			63556: outdata = 32'd1980;
			63557: outdata = 32'd1979;
			63558: outdata = 32'd1978;
			63559: outdata = 32'd1977;
			63560: outdata = 32'd1976;
			63561: outdata = 32'd1975;
			63562: outdata = 32'd1974;
			63563: outdata = 32'd1973;
			63564: outdata = 32'd1972;
			63565: outdata = 32'd1971;
			63566: outdata = 32'd1970;
			63567: outdata = 32'd1969;
			63568: outdata = 32'd1968;
			63569: outdata = 32'd1967;
			63570: outdata = 32'd1966;
			63571: outdata = 32'd1965;
			63572: outdata = 32'd1964;
			63573: outdata = 32'd1963;
			63574: outdata = 32'd1962;
			63575: outdata = 32'd1961;
			63576: outdata = 32'd1960;
			63577: outdata = 32'd1959;
			63578: outdata = 32'd1958;
			63579: outdata = 32'd1957;
			63580: outdata = 32'd1956;
			63581: outdata = 32'd1955;
			63582: outdata = 32'd1954;
			63583: outdata = 32'd1953;
			63584: outdata = 32'd1952;
			63585: outdata = 32'd1951;
			63586: outdata = 32'd1950;
			63587: outdata = 32'd1949;
			63588: outdata = 32'd1948;
			63589: outdata = 32'd1947;
			63590: outdata = 32'd1946;
			63591: outdata = 32'd1945;
			63592: outdata = 32'd1944;
			63593: outdata = 32'd1943;
			63594: outdata = 32'd1942;
			63595: outdata = 32'd1941;
			63596: outdata = 32'd1940;
			63597: outdata = 32'd1939;
			63598: outdata = 32'd1938;
			63599: outdata = 32'd1937;
			63600: outdata = 32'd1936;
			63601: outdata = 32'd1935;
			63602: outdata = 32'd1934;
			63603: outdata = 32'd1933;
			63604: outdata = 32'd1932;
			63605: outdata = 32'd1931;
			63606: outdata = 32'd1930;
			63607: outdata = 32'd1929;
			63608: outdata = 32'd1928;
			63609: outdata = 32'd1927;
			63610: outdata = 32'd1926;
			63611: outdata = 32'd1925;
			63612: outdata = 32'd1924;
			63613: outdata = 32'd1923;
			63614: outdata = 32'd1922;
			63615: outdata = 32'd1921;
			63616: outdata = 32'd1920;
			63617: outdata = 32'd1919;
			63618: outdata = 32'd1918;
			63619: outdata = 32'd1917;
			63620: outdata = 32'd1916;
			63621: outdata = 32'd1915;
			63622: outdata = 32'd1914;
			63623: outdata = 32'd1913;
			63624: outdata = 32'd1912;
			63625: outdata = 32'd1911;
			63626: outdata = 32'd1910;
			63627: outdata = 32'd1909;
			63628: outdata = 32'd1908;
			63629: outdata = 32'd1907;
			63630: outdata = 32'd1906;
			63631: outdata = 32'd1905;
			63632: outdata = 32'd1904;
			63633: outdata = 32'd1903;
			63634: outdata = 32'd1902;
			63635: outdata = 32'd1901;
			63636: outdata = 32'd1900;
			63637: outdata = 32'd1899;
			63638: outdata = 32'd1898;
			63639: outdata = 32'd1897;
			63640: outdata = 32'd1896;
			63641: outdata = 32'd1895;
			63642: outdata = 32'd1894;
			63643: outdata = 32'd1893;
			63644: outdata = 32'd1892;
			63645: outdata = 32'd1891;
			63646: outdata = 32'd1890;
			63647: outdata = 32'd1889;
			63648: outdata = 32'd1888;
			63649: outdata = 32'd1887;
			63650: outdata = 32'd1886;
			63651: outdata = 32'd1885;
			63652: outdata = 32'd1884;
			63653: outdata = 32'd1883;
			63654: outdata = 32'd1882;
			63655: outdata = 32'd1881;
			63656: outdata = 32'd1880;
			63657: outdata = 32'd1879;
			63658: outdata = 32'd1878;
			63659: outdata = 32'd1877;
			63660: outdata = 32'd1876;
			63661: outdata = 32'd1875;
			63662: outdata = 32'd1874;
			63663: outdata = 32'd1873;
			63664: outdata = 32'd1872;
			63665: outdata = 32'd1871;
			63666: outdata = 32'd1870;
			63667: outdata = 32'd1869;
			63668: outdata = 32'd1868;
			63669: outdata = 32'd1867;
			63670: outdata = 32'd1866;
			63671: outdata = 32'd1865;
			63672: outdata = 32'd1864;
			63673: outdata = 32'd1863;
			63674: outdata = 32'd1862;
			63675: outdata = 32'd1861;
			63676: outdata = 32'd1860;
			63677: outdata = 32'd1859;
			63678: outdata = 32'd1858;
			63679: outdata = 32'd1857;
			63680: outdata = 32'd1856;
			63681: outdata = 32'd1855;
			63682: outdata = 32'd1854;
			63683: outdata = 32'd1853;
			63684: outdata = 32'd1852;
			63685: outdata = 32'd1851;
			63686: outdata = 32'd1850;
			63687: outdata = 32'd1849;
			63688: outdata = 32'd1848;
			63689: outdata = 32'd1847;
			63690: outdata = 32'd1846;
			63691: outdata = 32'd1845;
			63692: outdata = 32'd1844;
			63693: outdata = 32'd1843;
			63694: outdata = 32'd1842;
			63695: outdata = 32'd1841;
			63696: outdata = 32'd1840;
			63697: outdata = 32'd1839;
			63698: outdata = 32'd1838;
			63699: outdata = 32'd1837;
			63700: outdata = 32'd1836;
			63701: outdata = 32'd1835;
			63702: outdata = 32'd1834;
			63703: outdata = 32'd1833;
			63704: outdata = 32'd1832;
			63705: outdata = 32'd1831;
			63706: outdata = 32'd1830;
			63707: outdata = 32'd1829;
			63708: outdata = 32'd1828;
			63709: outdata = 32'd1827;
			63710: outdata = 32'd1826;
			63711: outdata = 32'd1825;
			63712: outdata = 32'd1824;
			63713: outdata = 32'd1823;
			63714: outdata = 32'd1822;
			63715: outdata = 32'd1821;
			63716: outdata = 32'd1820;
			63717: outdata = 32'd1819;
			63718: outdata = 32'd1818;
			63719: outdata = 32'd1817;
			63720: outdata = 32'd1816;
			63721: outdata = 32'd1815;
			63722: outdata = 32'd1814;
			63723: outdata = 32'd1813;
			63724: outdata = 32'd1812;
			63725: outdata = 32'd1811;
			63726: outdata = 32'd1810;
			63727: outdata = 32'd1809;
			63728: outdata = 32'd1808;
			63729: outdata = 32'd1807;
			63730: outdata = 32'd1806;
			63731: outdata = 32'd1805;
			63732: outdata = 32'd1804;
			63733: outdata = 32'd1803;
			63734: outdata = 32'd1802;
			63735: outdata = 32'd1801;
			63736: outdata = 32'd1800;
			63737: outdata = 32'd1799;
			63738: outdata = 32'd1798;
			63739: outdata = 32'd1797;
			63740: outdata = 32'd1796;
			63741: outdata = 32'd1795;
			63742: outdata = 32'd1794;
			63743: outdata = 32'd1793;
			63744: outdata = 32'd1792;
			63745: outdata = 32'd1791;
			63746: outdata = 32'd1790;
			63747: outdata = 32'd1789;
			63748: outdata = 32'd1788;
			63749: outdata = 32'd1787;
			63750: outdata = 32'd1786;
			63751: outdata = 32'd1785;
			63752: outdata = 32'd1784;
			63753: outdata = 32'd1783;
			63754: outdata = 32'd1782;
			63755: outdata = 32'd1781;
			63756: outdata = 32'd1780;
			63757: outdata = 32'd1779;
			63758: outdata = 32'd1778;
			63759: outdata = 32'd1777;
			63760: outdata = 32'd1776;
			63761: outdata = 32'd1775;
			63762: outdata = 32'd1774;
			63763: outdata = 32'd1773;
			63764: outdata = 32'd1772;
			63765: outdata = 32'd1771;
			63766: outdata = 32'd1770;
			63767: outdata = 32'd1769;
			63768: outdata = 32'd1768;
			63769: outdata = 32'd1767;
			63770: outdata = 32'd1766;
			63771: outdata = 32'd1765;
			63772: outdata = 32'd1764;
			63773: outdata = 32'd1763;
			63774: outdata = 32'd1762;
			63775: outdata = 32'd1761;
			63776: outdata = 32'd1760;
			63777: outdata = 32'd1759;
			63778: outdata = 32'd1758;
			63779: outdata = 32'd1757;
			63780: outdata = 32'd1756;
			63781: outdata = 32'd1755;
			63782: outdata = 32'd1754;
			63783: outdata = 32'd1753;
			63784: outdata = 32'd1752;
			63785: outdata = 32'd1751;
			63786: outdata = 32'd1750;
			63787: outdata = 32'd1749;
			63788: outdata = 32'd1748;
			63789: outdata = 32'd1747;
			63790: outdata = 32'd1746;
			63791: outdata = 32'd1745;
			63792: outdata = 32'd1744;
			63793: outdata = 32'd1743;
			63794: outdata = 32'd1742;
			63795: outdata = 32'd1741;
			63796: outdata = 32'd1740;
			63797: outdata = 32'd1739;
			63798: outdata = 32'd1738;
			63799: outdata = 32'd1737;
			63800: outdata = 32'd1736;
			63801: outdata = 32'd1735;
			63802: outdata = 32'd1734;
			63803: outdata = 32'd1733;
			63804: outdata = 32'd1732;
			63805: outdata = 32'd1731;
			63806: outdata = 32'd1730;
			63807: outdata = 32'd1729;
			63808: outdata = 32'd1728;
			63809: outdata = 32'd1727;
			63810: outdata = 32'd1726;
			63811: outdata = 32'd1725;
			63812: outdata = 32'd1724;
			63813: outdata = 32'd1723;
			63814: outdata = 32'd1722;
			63815: outdata = 32'd1721;
			63816: outdata = 32'd1720;
			63817: outdata = 32'd1719;
			63818: outdata = 32'd1718;
			63819: outdata = 32'd1717;
			63820: outdata = 32'd1716;
			63821: outdata = 32'd1715;
			63822: outdata = 32'd1714;
			63823: outdata = 32'd1713;
			63824: outdata = 32'd1712;
			63825: outdata = 32'd1711;
			63826: outdata = 32'd1710;
			63827: outdata = 32'd1709;
			63828: outdata = 32'd1708;
			63829: outdata = 32'd1707;
			63830: outdata = 32'd1706;
			63831: outdata = 32'd1705;
			63832: outdata = 32'd1704;
			63833: outdata = 32'd1703;
			63834: outdata = 32'd1702;
			63835: outdata = 32'd1701;
			63836: outdata = 32'd1700;
			63837: outdata = 32'd1699;
			63838: outdata = 32'd1698;
			63839: outdata = 32'd1697;
			63840: outdata = 32'd1696;
			63841: outdata = 32'd1695;
			63842: outdata = 32'd1694;
			63843: outdata = 32'd1693;
			63844: outdata = 32'd1692;
			63845: outdata = 32'd1691;
			63846: outdata = 32'd1690;
			63847: outdata = 32'd1689;
			63848: outdata = 32'd1688;
			63849: outdata = 32'd1687;
			63850: outdata = 32'd1686;
			63851: outdata = 32'd1685;
			63852: outdata = 32'd1684;
			63853: outdata = 32'd1683;
			63854: outdata = 32'd1682;
			63855: outdata = 32'd1681;
			63856: outdata = 32'd1680;
			63857: outdata = 32'd1679;
			63858: outdata = 32'd1678;
			63859: outdata = 32'd1677;
			63860: outdata = 32'd1676;
			63861: outdata = 32'd1675;
			63862: outdata = 32'd1674;
			63863: outdata = 32'd1673;
			63864: outdata = 32'd1672;
			63865: outdata = 32'd1671;
			63866: outdata = 32'd1670;
			63867: outdata = 32'd1669;
			63868: outdata = 32'd1668;
			63869: outdata = 32'd1667;
			63870: outdata = 32'd1666;
			63871: outdata = 32'd1665;
			63872: outdata = 32'd1664;
			63873: outdata = 32'd1663;
			63874: outdata = 32'd1662;
			63875: outdata = 32'd1661;
			63876: outdata = 32'd1660;
			63877: outdata = 32'd1659;
			63878: outdata = 32'd1658;
			63879: outdata = 32'd1657;
			63880: outdata = 32'd1656;
			63881: outdata = 32'd1655;
			63882: outdata = 32'd1654;
			63883: outdata = 32'd1653;
			63884: outdata = 32'd1652;
			63885: outdata = 32'd1651;
			63886: outdata = 32'd1650;
			63887: outdata = 32'd1649;
			63888: outdata = 32'd1648;
			63889: outdata = 32'd1647;
			63890: outdata = 32'd1646;
			63891: outdata = 32'd1645;
			63892: outdata = 32'd1644;
			63893: outdata = 32'd1643;
			63894: outdata = 32'd1642;
			63895: outdata = 32'd1641;
			63896: outdata = 32'd1640;
			63897: outdata = 32'd1639;
			63898: outdata = 32'd1638;
			63899: outdata = 32'd1637;
			63900: outdata = 32'd1636;
			63901: outdata = 32'd1635;
			63902: outdata = 32'd1634;
			63903: outdata = 32'd1633;
			63904: outdata = 32'd1632;
			63905: outdata = 32'd1631;
			63906: outdata = 32'd1630;
			63907: outdata = 32'd1629;
			63908: outdata = 32'd1628;
			63909: outdata = 32'd1627;
			63910: outdata = 32'd1626;
			63911: outdata = 32'd1625;
			63912: outdata = 32'd1624;
			63913: outdata = 32'd1623;
			63914: outdata = 32'd1622;
			63915: outdata = 32'd1621;
			63916: outdata = 32'd1620;
			63917: outdata = 32'd1619;
			63918: outdata = 32'd1618;
			63919: outdata = 32'd1617;
			63920: outdata = 32'd1616;
			63921: outdata = 32'd1615;
			63922: outdata = 32'd1614;
			63923: outdata = 32'd1613;
			63924: outdata = 32'd1612;
			63925: outdata = 32'd1611;
			63926: outdata = 32'd1610;
			63927: outdata = 32'd1609;
			63928: outdata = 32'd1608;
			63929: outdata = 32'd1607;
			63930: outdata = 32'd1606;
			63931: outdata = 32'd1605;
			63932: outdata = 32'd1604;
			63933: outdata = 32'd1603;
			63934: outdata = 32'd1602;
			63935: outdata = 32'd1601;
			63936: outdata = 32'd1600;
			63937: outdata = 32'd1599;
			63938: outdata = 32'd1598;
			63939: outdata = 32'd1597;
			63940: outdata = 32'd1596;
			63941: outdata = 32'd1595;
			63942: outdata = 32'd1594;
			63943: outdata = 32'd1593;
			63944: outdata = 32'd1592;
			63945: outdata = 32'd1591;
			63946: outdata = 32'd1590;
			63947: outdata = 32'd1589;
			63948: outdata = 32'd1588;
			63949: outdata = 32'd1587;
			63950: outdata = 32'd1586;
			63951: outdata = 32'd1585;
			63952: outdata = 32'd1584;
			63953: outdata = 32'd1583;
			63954: outdata = 32'd1582;
			63955: outdata = 32'd1581;
			63956: outdata = 32'd1580;
			63957: outdata = 32'd1579;
			63958: outdata = 32'd1578;
			63959: outdata = 32'd1577;
			63960: outdata = 32'd1576;
			63961: outdata = 32'd1575;
			63962: outdata = 32'd1574;
			63963: outdata = 32'd1573;
			63964: outdata = 32'd1572;
			63965: outdata = 32'd1571;
			63966: outdata = 32'd1570;
			63967: outdata = 32'd1569;
			63968: outdata = 32'd1568;
			63969: outdata = 32'd1567;
			63970: outdata = 32'd1566;
			63971: outdata = 32'd1565;
			63972: outdata = 32'd1564;
			63973: outdata = 32'd1563;
			63974: outdata = 32'd1562;
			63975: outdata = 32'd1561;
			63976: outdata = 32'd1560;
			63977: outdata = 32'd1559;
			63978: outdata = 32'd1558;
			63979: outdata = 32'd1557;
			63980: outdata = 32'd1556;
			63981: outdata = 32'd1555;
			63982: outdata = 32'd1554;
			63983: outdata = 32'd1553;
			63984: outdata = 32'd1552;
			63985: outdata = 32'd1551;
			63986: outdata = 32'd1550;
			63987: outdata = 32'd1549;
			63988: outdata = 32'd1548;
			63989: outdata = 32'd1547;
			63990: outdata = 32'd1546;
			63991: outdata = 32'd1545;
			63992: outdata = 32'd1544;
			63993: outdata = 32'd1543;
			63994: outdata = 32'd1542;
			63995: outdata = 32'd1541;
			63996: outdata = 32'd1540;
			63997: outdata = 32'd1539;
			63998: outdata = 32'd1538;
			63999: outdata = 32'd1537;
			64000: outdata = 32'd1536;
			64001: outdata = 32'd1535;
			64002: outdata = 32'd1534;
			64003: outdata = 32'd1533;
			64004: outdata = 32'd1532;
			64005: outdata = 32'd1531;
			64006: outdata = 32'd1530;
			64007: outdata = 32'd1529;
			64008: outdata = 32'd1528;
			64009: outdata = 32'd1527;
			64010: outdata = 32'd1526;
			64011: outdata = 32'd1525;
			64012: outdata = 32'd1524;
			64013: outdata = 32'd1523;
			64014: outdata = 32'd1522;
			64015: outdata = 32'd1521;
			64016: outdata = 32'd1520;
			64017: outdata = 32'd1519;
			64018: outdata = 32'd1518;
			64019: outdata = 32'd1517;
			64020: outdata = 32'd1516;
			64021: outdata = 32'd1515;
			64022: outdata = 32'd1514;
			64023: outdata = 32'd1513;
			64024: outdata = 32'd1512;
			64025: outdata = 32'd1511;
			64026: outdata = 32'd1510;
			64027: outdata = 32'd1509;
			64028: outdata = 32'd1508;
			64029: outdata = 32'd1507;
			64030: outdata = 32'd1506;
			64031: outdata = 32'd1505;
			64032: outdata = 32'd1504;
			64033: outdata = 32'd1503;
			64034: outdata = 32'd1502;
			64035: outdata = 32'd1501;
			64036: outdata = 32'd1500;
			64037: outdata = 32'd1499;
			64038: outdata = 32'd1498;
			64039: outdata = 32'd1497;
			64040: outdata = 32'd1496;
			64041: outdata = 32'd1495;
			64042: outdata = 32'd1494;
			64043: outdata = 32'd1493;
			64044: outdata = 32'd1492;
			64045: outdata = 32'd1491;
			64046: outdata = 32'd1490;
			64047: outdata = 32'd1489;
			64048: outdata = 32'd1488;
			64049: outdata = 32'd1487;
			64050: outdata = 32'd1486;
			64051: outdata = 32'd1485;
			64052: outdata = 32'd1484;
			64053: outdata = 32'd1483;
			64054: outdata = 32'd1482;
			64055: outdata = 32'd1481;
			64056: outdata = 32'd1480;
			64057: outdata = 32'd1479;
			64058: outdata = 32'd1478;
			64059: outdata = 32'd1477;
			64060: outdata = 32'd1476;
			64061: outdata = 32'd1475;
			64062: outdata = 32'd1474;
			64063: outdata = 32'd1473;
			64064: outdata = 32'd1472;
			64065: outdata = 32'd1471;
			64066: outdata = 32'd1470;
			64067: outdata = 32'd1469;
			64068: outdata = 32'd1468;
			64069: outdata = 32'd1467;
			64070: outdata = 32'd1466;
			64071: outdata = 32'd1465;
			64072: outdata = 32'd1464;
			64073: outdata = 32'd1463;
			64074: outdata = 32'd1462;
			64075: outdata = 32'd1461;
			64076: outdata = 32'd1460;
			64077: outdata = 32'd1459;
			64078: outdata = 32'd1458;
			64079: outdata = 32'd1457;
			64080: outdata = 32'd1456;
			64081: outdata = 32'd1455;
			64082: outdata = 32'd1454;
			64083: outdata = 32'd1453;
			64084: outdata = 32'd1452;
			64085: outdata = 32'd1451;
			64086: outdata = 32'd1450;
			64087: outdata = 32'd1449;
			64088: outdata = 32'd1448;
			64089: outdata = 32'd1447;
			64090: outdata = 32'd1446;
			64091: outdata = 32'd1445;
			64092: outdata = 32'd1444;
			64093: outdata = 32'd1443;
			64094: outdata = 32'd1442;
			64095: outdata = 32'd1441;
			64096: outdata = 32'd1440;
			64097: outdata = 32'd1439;
			64098: outdata = 32'd1438;
			64099: outdata = 32'd1437;
			64100: outdata = 32'd1436;
			64101: outdata = 32'd1435;
			64102: outdata = 32'd1434;
			64103: outdata = 32'd1433;
			64104: outdata = 32'd1432;
			64105: outdata = 32'd1431;
			64106: outdata = 32'd1430;
			64107: outdata = 32'd1429;
			64108: outdata = 32'd1428;
			64109: outdata = 32'd1427;
			64110: outdata = 32'd1426;
			64111: outdata = 32'd1425;
			64112: outdata = 32'd1424;
			64113: outdata = 32'd1423;
			64114: outdata = 32'd1422;
			64115: outdata = 32'd1421;
			64116: outdata = 32'd1420;
			64117: outdata = 32'd1419;
			64118: outdata = 32'd1418;
			64119: outdata = 32'd1417;
			64120: outdata = 32'd1416;
			64121: outdata = 32'd1415;
			64122: outdata = 32'd1414;
			64123: outdata = 32'd1413;
			64124: outdata = 32'd1412;
			64125: outdata = 32'd1411;
			64126: outdata = 32'd1410;
			64127: outdata = 32'd1409;
			64128: outdata = 32'd1408;
			64129: outdata = 32'd1407;
			64130: outdata = 32'd1406;
			64131: outdata = 32'd1405;
			64132: outdata = 32'd1404;
			64133: outdata = 32'd1403;
			64134: outdata = 32'd1402;
			64135: outdata = 32'd1401;
			64136: outdata = 32'd1400;
			64137: outdata = 32'd1399;
			64138: outdata = 32'd1398;
			64139: outdata = 32'd1397;
			64140: outdata = 32'd1396;
			64141: outdata = 32'd1395;
			64142: outdata = 32'd1394;
			64143: outdata = 32'd1393;
			64144: outdata = 32'd1392;
			64145: outdata = 32'd1391;
			64146: outdata = 32'd1390;
			64147: outdata = 32'd1389;
			64148: outdata = 32'd1388;
			64149: outdata = 32'd1387;
			64150: outdata = 32'd1386;
			64151: outdata = 32'd1385;
			64152: outdata = 32'd1384;
			64153: outdata = 32'd1383;
			64154: outdata = 32'd1382;
			64155: outdata = 32'd1381;
			64156: outdata = 32'd1380;
			64157: outdata = 32'd1379;
			64158: outdata = 32'd1378;
			64159: outdata = 32'd1377;
			64160: outdata = 32'd1376;
			64161: outdata = 32'd1375;
			64162: outdata = 32'd1374;
			64163: outdata = 32'd1373;
			64164: outdata = 32'd1372;
			64165: outdata = 32'd1371;
			64166: outdata = 32'd1370;
			64167: outdata = 32'd1369;
			64168: outdata = 32'd1368;
			64169: outdata = 32'd1367;
			64170: outdata = 32'd1366;
			64171: outdata = 32'd1365;
			64172: outdata = 32'd1364;
			64173: outdata = 32'd1363;
			64174: outdata = 32'd1362;
			64175: outdata = 32'd1361;
			64176: outdata = 32'd1360;
			64177: outdata = 32'd1359;
			64178: outdata = 32'd1358;
			64179: outdata = 32'd1357;
			64180: outdata = 32'd1356;
			64181: outdata = 32'd1355;
			64182: outdata = 32'd1354;
			64183: outdata = 32'd1353;
			64184: outdata = 32'd1352;
			64185: outdata = 32'd1351;
			64186: outdata = 32'd1350;
			64187: outdata = 32'd1349;
			64188: outdata = 32'd1348;
			64189: outdata = 32'd1347;
			64190: outdata = 32'd1346;
			64191: outdata = 32'd1345;
			64192: outdata = 32'd1344;
			64193: outdata = 32'd1343;
			64194: outdata = 32'd1342;
			64195: outdata = 32'd1341;
			64196: outdata = 32'd1340;
			64197: outdata = 32'd1339;
			64198: outdata = 32'd1338;
			64199: outdata = 32'd1337;
			64200: outdata = 32'd1336;
			64201: outdata = 32'd1335;
			64202: outdata = 32'd1334;
			64203: outdata = 32'd1333;
			64204: outdata = 32'd1332;
			64205: outdata = 32'd1331;
			64206: outdata = 32'd1330;
			64207: outdata = 32'd1329;
			64208: outdata = 32'd1328;
			64209: outdata = 32'd1327;
			64210: outdata = 32'd1326;
			64211: outdata = 32'd1325;
			64212: outdata = 32'd1324;
			64213: outdata = 32'd1323;
			64214: outdata = 32'd1322;
			64215: outdata = 32'd1321;
			64216: outdata = 32'd1320;
			64217: outdata = 32'd1319;
			64218: outdata = 32'd1318;
			64219: outdata = 32'd1317;
			64220: outdata = 32'd1316;
			64221: outdata = 32'd1315;
			64222: outdata = 32'd1314;
			64223: outdata = 32'd1313;
			64224: outdata = 32'd1312;
			64225: outdata = 32'd1311;
			64226: outdata = 32'd1310;
			64227: outdata = 32'd1309;
			64228: outdata = 32'd1308;
			64229: outdata = 32'd1307;
			64230: outdata = 32'd1306;
			64231: outdata = 32'd1305;
			64232: outdata = 32'd1304;
			64233: outdata = 32'd1303;
			64234: outdata = 32'd1302;
			64235: outdata = 32'd1301;
			64236: outdata = 32'd1300;
			64237: outdata = 32'd1299;
			64238: outdata = 32'd1298;
			64239: outdata = 32'd1297;
			64240: outdata = 32'd1296;
			64241: outdata = 32'd1295;
			64242: outdata = 32'd1294;
			64243: outdata = 32'd1293;
			64244: outdata = 32'd1292;
			64245: outdata = 32'd1291;
			64246: outdata = 32'd1290;
			64247: outdata = 32'd1289;
			64248: outdata = 32'd1288;
			64249: outdata = 32'd1287;
			64250: outdata = 32'd1286;
			64251: outdata = 32'd1285;
			64252: outdata = 32'd1284;
			64253: outdata = 32'd1283;
			64254: outdata = 32'd1282;
			64255: outdata = 32'd1281;
			64256: outdata = 32'd1280;
			64257: outdata = 32'd1279;
			64258: outdata = 32'd1278;
			64259: outdata = 32'd1277;
			64260: outdata = 32'd1276;
			64261: outdata = 32'd1275;
			64262: outdata = 32'd1274;
			64263: outdata = 32'd1273;
			64264: outdata = 32'd1272;
			64265: outdata = 32'd1271;
			64266: outdata = 32'd1270;
			64267: outdata = 32'd1269;
			64268: outdata = 32'd1268;
			64269: outdata = 32'd1267;
			64270: outdata = 32'd1266;
			64271: outdata = 32'd1265;
			64272: outdata = 32'd1264;
			64273: outdata = 32'd1263;
			64274: outdata = 32'd1262;
			64275: outdata = 32'd1261;
			64276: outdata = 32'd1260;
			64277: outdata = 32'd1259;
			64278: outdata = 32'd1258;
			64279: outdata = 32'd1257;
			64280: outdata = 32'd1256;
			64281: outdata = 32'd1255;
			64282: outdata = 32'd1254;
			64283: outdata = 32'd1253;
			64284: outdata = 32'd1252;
			64285: outdata = 32'd1251;
			64286: outdata = 32'd1250;
			64287: outdata = 32'd1249;
			64288: outdata = 32'd1248;
			64289: outdata = 32'd1247;
			64290: outdata = 32'd1246;
			64291: outdata = 32'd1245;
			64292: outdata = 32'd1244;
			64293: outdata = 32'd1243;
			64294: outdata = 32'd1242;
			64295: outdata = 32'd1241;
			64296: outdata = 32'd1240;
			64297: outdata = 32'd1239;
			64298: outdata = 32'd1238;
			64299: outdata = 32'd1237;
			64300: outdata = 32'd1236;
			64301: outdata = 32'd1235;
			64302: outdata = 32'd1234;
			64303: outdata = 32'd1233;
			64304: outdata = 32'd1232;
			64305: outdata = 32'd1231;
			64306: outdata = 32'd1230;
			64307: outdata = 32'd1229;
			64308: outdata = 32'd1228;
			64309: outdata = 32'd1227;
			64310: outdata = 32'd1226;
			64311: outdata = 32'd1225;
			64312: outdata = 32'd1224;
			64313: outdata = 32'd1223;
			64314: outdata = 32'd1222;
			64315: outdata = 32'd1221;
			64316: outdata = 32'd1220;
			64317: outdata = 32'd1219;
			64318: outdata = 32'd1218;
			64319: outdata = 32'd1217;
			64320: outdata = 32'd1216;
			64321: outdata = 32'd1215;
			64322: outdata = 32'd1214;
			64323: outdata = 32'd1213;
			64324: outdata = 32'd1212;
			64325: outdata = 32'd1211;
			64326: outdata = 32'd1210;
			64327: outdata = 32'd1209;
			64328: outdata = 32'd1208;
			64329: outdata = 32'd1207;
			64330: outdata = 32'd1206;
			64331: outdata = 32'd1205;
			64332: outdata = 32'd1204;
			64333: outdata = 32'd1203;
			64334: outdata = 32'd1202;
			64335: outdata = 32'd1201;
			64336: outdata = 32'd1200;
			64337: outdata = 32'd1199;
			64338: outdata = 32'd1198;
			64339: outdata = 32'd1197;
			64340: outdata = 32'd1196;
			64341: outdata = 32'd1195;
			64342: outdata = 32'd1194;
			64343: outdata = 32'd1193;
			64344: outdata = 32'd1192;
			64345: outdata = 32'd1191;
			64346: outdata = 32'd1190;
			64347: outdata = 32'd1189;
			64348: outdata = 32'd1188;
			64349: outdata = 32'd1187;
			64350: outdata = 32'd1186;
			64351: outdata = 32'd1185;
			64352: outdata = 32'd1184;
			64353: outdata = 32'd1183;
			64354: outdata = 32'd1182;
			64355: outdata = 32'd1181;
			64356: outdata = 32'd1180;
			64357: outdata = 32'd1179;
			64358: outdata = 32'd1178;
			64359: outdata = 32'd1177;
			64360: outdata = 32'd1176;
			64361: outdata = 32'd1175;
			64362: outdata = 32'd1174;
			64363: outdata = 32'd1173;
			64364: outdata = 32'd1172;
			64365: outdata = 32'd1171;
			64366: outdata = 32'd1170;
			64367: outdata = 32'd1169;
			64368: outdata = 32'd1168;
			64369: outdata = 32'd1167;
			64370: outdata = 32'd1166;
			64371: outdata = 32'd1165;
			64372: outdata = 32'd1164;
			64373: outdata = 32'd1163;
			64374: outdata = 32'd1162;
			64375: outdata = 32'd1161;
			64376: outdata = 32'd1160;
			64377: outdata = 32'd1159;
			64378: outdata = 32'd1158;
			64379: outdata = 32'd1157;
			64380: outdata = 32'd1156;
			64381: outdata = 32'd1155;
			64382: outdata = 32'd1154;
			64383: outdata = 32'd1153;
			64384: outdata = 32'd1152;
			64385: outdata = 32'd1151;
			64386: outdata = 32'd1150;
			64387: outdata = 32'd1149;
			64388: outdata = 32'd1148;
			64389: outdata = 32'd1147;
			64390: outdata = 32'd1146;
			64391: outdata = 32'd1145;
			64392: outdata = 32'd1144;
			64393: outdata = 32'd1143;
			64394: outdata = 32'd1142;
			64395: outdata = 32'd1141;
			64396: outdata = 32'd1140;
			64397: outdata = 32'd1139;
			64398: outdata = 32'd1138;
			64399: outdata = 32'd1137;
			64400: outdata = 32'd1136;
			64401: outdata = 32'd1135;
			64402: outdata = 32'd1134;
			64403: outdata = 32'd1133;
			64404: outdata = 32'd1132;
			64405: outdata = 32'd1131;
			64406: outdata = 32'd1130;
			64407: outdata = 32'd1129;
			64408: outdata = 32'd1128;
			64409: outdata = 32'd1127;
			64410: outdata = 32'd1126;
			64411: outdata = 32'd1125;
			64412: outdata = 32'd1124;
			64413: outdata = 32'd1123;
			64414: outdata = 32'd1122;
			64415: outdata = 32'd1121;
			64416: outdata = 32'd1120;
			64417: outdata = 32'd1119;
			64418: outdata = 32'd1118;
			64419: outdata = 32'd1117;
			64420: outdata = 32'd1116;
			64421: outdata = 32'd1115;
			64422: outdata = 32'd1114;
			64423: outdata = 32'd1113;
			64424: outdata = 32'd1112;
			64425: outdata = 32'd1111;
			64426: outdata = 32'd1110;
			64427: outdata = 32'd1109;
			64428: outdata = 32'd1108;
			64429: outdata = 32'd1107;
			64430: outdata = 32'd1106;
			64431: outdata = 32'd1105;
			64432: outdata = 32'd1104;
			64433: outdata = 32'd1103;
			64434: outdata = 32'd1102;
			64435: outdata = 32'd1101;
			64436: outdata = 32'd1100;
			64437: outdata = 32'd1099;
			64438: outdata = 32'd1098;
			64439: outdata = 32'd1097;
			64440: outdata = 32'd1096;
			64441: outdata = 32'd1095;
			64442: outdata = 32'd1094;
			64443: outdata = 32'd1093;
			64444: outdata = 32'd1092;
			64445: outdata = 32'd1091;
			64446: outdata = 32'd1090;
			64447: outdata = 32'd1089;
			64448: outdata = 32'd1088;
			64449: outdata = 32'd1087;
			64450: outdata = 32'd1086;
			64451: outdata = 32'd1085;
			64452: outdata = 32'd1084;
			64453: outdata = 32'd1083;
			64454: outdata = 32'd1082;
			64455: outdata = 32'd1081;
			64456: outdata = 32'd1080;
			64457: outdata = 32'd1079;
			64458: outdata = 32'd1078;
			64459: outdata = 32'd1077;
			64460: outdata = 32'd1076;
			64461: outdata = 32'd1075;
			64462: outdata = 32'd1074;
			64463: outdata = 32'd1073;
			64464: outdata = 32'd1072;
			64465: outdata = 32'd1071;
			64466: outdata = 32'd1070;
			64467: outdata = 32'd1069;
			64468: outdata = 32'd1068;
			64469: outdata = 32'd1067;
			64470: outdata = 32'd1066;
			64471: outdata = 32'd1065;
			64472: outdata = 32'd1064;
			64473: outdata = 32'd1063;
			64474: outdata = 32'd1062;
			64475: outdata = 32'd1061;
			64476: outdata = 32'd1060;
			64477: outdata = 32'd1059;
			64478: outdata = 32'd1058;
			64479: outdata = 32'd1057;
			64480: outdata = 32'd1056;
			64481: outdata = 32'd1055;
			64482: outdata = 32'd1054;
			64483: outdata = 32'd1053;
			64484: outdata = 32'd1052;
			64485: outdata = 32'd1051;
			64486: outdata = 32'd1050;
			64487: outdata = 32'd1049;
			64488: outdata = 32'd1048;
			64489: outdata = 32'd1047;
			64490: outdata = 32'd1046;
			64491: outdata = 32'd1045;
			64492: outdata = 32'd1044;
			64493: outdata = 32'd1043;
			64494: outdata = 32'd1042;
			64495: outdata = 32'd1041;
			64496: outdata = 32'd1040;
			64497: outdata = 32'd1039;
			64498: outdata = 32'd1038;
			64499: outdata = 32'd1037;
			64500: outdata = 32'd1036;
			64501: outdata = 32'd1035;
			64502: outdata = 32'd1034;
			64503: outdata = 32'd1033;
			64504: outdata = 32'd1032;
			64505: outdata = 32'd1031;
			64506: outdata = 32'd1030;
			64507: outdata = 32'd1029;
			64508: outdata = 32'd1028;
			64509: outdata = 32'd1027;
			64510: outdata = 32'd1026;
			64511: outdata = 32'd1025;
			64512: outdata = 32'd1024;
			64513: outdata = 32'd1023;
			64514: outdata = 32'd1022;
			64515: outdata = 32'd1021;
			64516: outdata = 32'd1020;
			64517: outdata = 32'd1019;
			64518: outdata = 32'd1018;
			64519: outdata = 32'd1017;
			64520: outdata = 32'd1016;
			64521: outdata = 32'd1015;
			64522: outdata = 32'd1014;
			64523: outdata = 32'd1013;
			64524: outdata = 32'd1012;
			64525: outdata = 32'd1011;
			64526: outdata = 32'd1010;
			64527: outdata = 32'd1009;
			64528: outdata = 32'd1008;
			64529: outdata = 32'd1007;
			64530: outdata = 32'd1006;
			64531: outdata = 32'd1005;
			64532: outdata = 32'd1004;
			64533: outdata = 32'd1003;
			64534: outdata = 32'd1002;
			64535: outdata = 32'd1001;
			64536: outdata = 32'd1000;
			64537: outdata = 32'd999;
			64538: outdata = 32'd998;
			64539: outdata = 32'd997;
			64540: outdata = 32'd996;
			64541: outdata = 32'd995;
			64542: outdata = 32'd994;
			64543: outdata = 32'd993;
			64544: outdata = 32'd992;
			64545: outdata = 32'd991;
			64546: outdata = 32'd990;
			64547: outdata = 32'd989;
			64548: outdata = 32'd988;
			64549: outdata = 32'd987;
			64550: outdata = 32'd986;
			64551: outdata = 32'd985;
			64552: outdata = 32'd984;
			64553: outdata = 32'd983;
			64554: outdata = 32'd982;
			64555: outdata = 32'd981;
			64556: outdata = 32'd980;
			64557: outdata = 32'd979;
			64558: outdata = 32'd978;
			64559: outdata = 32'd977;
			64560: outdata = 32'd976;
			64561: outdata = 32'd975;
			64562: outdata = 32'd974;
			64563: outdata = 32'd973;
			64564: outdata = 32'd972;
			64565: outdata = 32'd971;
			64566: outdata = 32'd970;
			64567: outdata = 32'd969;
			64568: outdata = 32'd968;
			64569: outdata = 32'd967;
			64570: outdata = 32'd966;
			64571: outdata = 32'd965;
			64572: outdata = 32'd964;
			64573: outdata = 32'd963;
			64574: outdata = 32'd962;
			64575: outdata = 32'd961;
			64576: outdata = 32'd960;
			64577: outdata = 32'd959;
			64578: outdata = 32'd958;
			64579: outdata = 32'd957;
			64580: outdata = 32'd956;
			64581: outdata = 32'd955;
			64582: outdata = 32'd954;
			64583: outdata = 32'd953;
			64584: outdata = 32'd952;
			64585: outdata = 32'd951;
			64586: outdata = 32'd950;
			64587: outdata = 32'd949;
			64588: outdata = 32'd948;
			64589: outdata = 32'd947;
			64590: outdata = 32'd946;
			64591: outdata = 32'd945;
			64592: outdata = 32'd944;
			64593: outdata = 32'd943;
			64594: outdata = 32'd942;
			64595: outdata = 32'd941;
			64596: outdata = 32'd940;
			64597: outdata = 32'd939;
			64598: outdata = 32'd938;
			64599: outdata = 32'd937;
			64600: outdata = 32'd936;
			64601: outdata = 32'd935;
			64602: outdata = 32'd934;
			64603: outdata = 32'd933;
			64604: outdata = 32'd932;
			64605: outdata = 32'd931;
			64606: outdata = 32'd930;
			64607: outdata = 32'd929;
			64608: outdata = 32'd928;
			64609: outdata = 32'd927;
			64610: outdata = 32'd926;
			64611: outdata = 32'd925;
			64612: outdata = 32'd924;
			64613: outdata = 32'd923;
			64614: outdata = 32'd922;
			64615: outdata = 32'd921;
			64616: outdata = 32'd920;
			64617: outdata = 32'd919;
			64618: outdata = 32'd918;
			64619: outdata = 32'd917;
			64620: outdata = 32'd916;
			64621: outdata = 32'd915;
			64622: outdata = 32'd914;
			64623: outdata = 32'd913;
			64624: outdata = 32'd912;
			64625: outdata = 32'd911;
			64626: outdata = 32'd910;
			64627: outdata = 32'd909;
			64628: outdata = 32'd908;
			64629: outdata = 32'd907;
			64630: outdata = 32'd906;
			64631: outdata = 32'd905;
			64632: outdata = 32'd904;
			64633: outdata = 32'd903;
			64634: outdata = 32'd902;
			64635: outdata = 32'd901;
			64636: outdata = 32'd900;
			64637: outdata = 32'd899;
			64638: outdata = 32'd898;
			64639: outdata = 32'd897;
			64640: outdata = 32'd896;
			64641: outdata = 32'd895;
			64642: outdata = 32'd894;
			64643: outdata = 32'd893;
			64644: outdata = 32'd892;
			64645: outdata = 32'd891;
			64646: outdata = 32'd890;
			64647: outdata = 32'd889;
			64648: outdata = 32'd888;
			64649: outdata = 32'd887;
			64650: outdata = 32'd886;
			64651: outdata = 32'd885;
			64652: outdata = 32'd884;
			64653: outdata = 32'd883;
			64654: outdata = 32'd882;
			64655: outdata = 32'd881;
			64656: outdata = 32'd880;
			64657: outdata = 32'd879;
			64658: outdata = 32'd878;
			64659: outdata = 32'd877;
			64660: outdata = 32'd876;
			64661: outdata = 32'd875;
			64662: outdata = 32'd874;
			64663: outdata = 32'd873;
			64664: outdata = 32'd872;
			64665: outdata = 32'd871;
			64666: outdata = 32'd870;
			64667: outdata = 32'd869;
			64668: outdata = 32'd868;
			64669: outdata = 32'd867;
			64670: outdata = 32'd866;
			64671: outdata = 32'd865;
			64672: outdata = 32'd864;
			64673: outdata = 32'd863;
			64674: outdata = 32'd862;
			64675: outdata = 32'd861;
			64676: outdata = 32'd860;
			64677: outdata = 32'd859;
			64678: outdata = 32'd858;
			64679: outdata = 32'd857;
			64680: outdata = 32'd856;
			64681: outdata = 32'd855;
			64682: outdata = 32'd854;
			64683: outdata = 32'd853;
			64684: outdata = 32'd852;
			64685: outdata = 32'd851;
			64686: outdata = 32'd850;
			64687: outdata = 32'd849;
			64688: outdata = 32'd848;
			64689: outdata = 32'd847;
			64690: outdata = 32'd846;
			64691: outdata = 32'd845;
			64692: outdata = 32'd844;
			64693: outdata = 32'd843;
			64694: outdata = 32'd842;
			64695: outdata = 32'd841;
			64696: outdata = 32'd840;
			64697: outdata = 32'd839;
			64698: outdata = 32'd838;
			64699: outdata = 32'd837;
			64700: outdata = 32'd836;
			64701: outdata = 32'd835;
			64702: outdata = 32'd834;
			64703: outdata = 32'd833;
			64704: outdata = 32'd832;
			64705: outdata = 32'd831;
			64706: outdata = 32'd830;
			64707: outdata = 32'd829;
			64708: outdata = 32'd828;
			64709: outdata = 32'd827;
			64710: outdata = 32'd826;
			64711: outdata = 32'd825;
			64712: outdata = 32'd824;
			64713: outdata = 32'd823;
			64714: outdata = 32'd822;
			64715: outdata = 32'd821;
			64716: outdata = 32'd820;
			64717: outdata = 32'd819;
			64718: outdata = 32'd818;
			64719: outdata = 32'd817;
			64720: outdata = 32'd816;
			64721: outdata = 32'd815;
			64722: outdata = 32'd814;
			64723: outdata = 32'd813;
			64724: outdata = 32'd812;
			64725: outdata = 32'd811;
			64726: outdata = 32'd810;
			64727: outdata = 32'd809;
			64728: outdata = 32'd808;
			64729: outdata = 32'd807;
			64730: outdata = 32'd806;
			64731: outdata = 32'd805;
			64732: outdata = 32'd804;
			64733: outdata = 32'd803;
			64734: outdata = 32'd802;
			64735: outdata = 32'd801;
			64736: outdata = 32'd800;
			64737: outdata = 32'd799;
			64738: outdata = 32'd798;
			64739: outdata = 32'd797;
			64740: outdata = 32'd796;
			64741: outdata = 32'd795;
			64742: outdata = 32'd794;
			64743: outdata = 32'd793;
			64744: outdata = 32'd792;
			64745: outdata = 32'd791;
			64746: outdata = 32'd790;
			64747: outdata = 32'd789;
			64748: outdata = 32'd788;
			64749: outdata = 32'd787;
			64750: outdata = 32'd786;
			64751: outdata = 32'd785;
			64752: outdata = 32'd784;
			64753: outdata = 32'd783;
			64754: outdata = 32'd782;
			64755: outdata = 32'd781;
			64756: outdata = 32'd780;
			64757: outdata = 32'd779;
			64758: outdata = 32'd778;
			64759: outdata = 32'd777;
			64760: outdata = 32'd776;
			64761: outdata = 32'd775;
			64762: outdata = 32'd774;
			64763: outdata = 32'd773;
			64764: outdata = 32'd772;
			64765: outdata = 32'd771;
			64766: outdata = 32'd770;
			64767: outdata = 32'd769;
			64768: outdata = 32'd768;
			64769: outdata = 32'd767;
			64770: outdata = 32'd766;
			64771: outdata = 32'd765;
			64772: outdata = 32'd764;
			64773: outdata = 32'd763;
			64774: outdata = 32'd762;
			64775: outdata = 32'd761;
			64776: outdata = 32'd760;
			64777: outdata = 32'd759;
			64778: outdata = 32'd758;
			64779: outdata = 32'd757;
			64780: outdata = 32'd756;
			64781: outdata = 32'd755;
			64782: outdata = 32'd754;
			64783: outdata = 32'd753;
			64784: outdata = 32'd752;
			64785: outdata = 32'd751;
			64786: outdata = 32'd750;
			64787: outdata = 32'd749;
			64788: outdata = 32'd748;
			64789: outdata = 32'd747;
			64790: outdata = 32'd746;
			64791: outdata = 32'd745;
			64792: outdata = 32'd744;
			64793: outdata = 32'd743;
			64794: outdata = 32'd742;
			64795: outdata = 32'd741;
			64796: outdata = 32'd740;
			64797: outdata = 32'd739;
			64798: outdata = 32'd738;
			64799: outdata = 32'd737;
			64800: outdata = 32'd736;
			64801: outdata = 32'd735;
			64802: outdata = 32'd734;
			64803: outdata = 32'd733;
			64804: outdata = 32'd732;
			64805: outdata = 32'd731;
			64806: outdata = 32'd730;
			64807: outdata = 32'd729;
			64808: outdata = 32'd728;
			64809: outdata = 32'd727;
			64810: outdata = 32'd726;
			64811: outdata = 32'd725;
			64812: outdata = 32'd724;
			64813: outdata = 32'd723;
			64814: outdata = 32'd722;
			64815: outdata = 32'd721;
			64816: outdata = 32'd720;
			64817: outdata = 32'd719;
			64818: outdata = 32'd718;
			64819: outdata = 32'd717;
			64820: outdata = 32'd716;
			64821: outdata = 32'd715;
			64822: outdata = 32'd714;
			64823: outdata = 32'd713;
			64824: outdata = 32'd712;
			64825: outdata = 32'd711;
			64826: outdata = 32'd710;
			64827: outdata = 32'd709;
			64828: outdata = 32'd708;
			64829: outdata = 32'd707;
			64830: outdata = 32'd706;
			64831: outdata = 32'd705;
			64832: outdata = 32'd704;
			64833: outdata = 32'd703;
			64834: outdata = 32'd702;
			64835: outdata = 32'd701;
			64836: outdata = 32'd700;
			64837: outdata = 32'd699;
			64838: outdata = 32'd698;
			64839: outdata = 32'd697;
			64840: outdata = 32'd696;
			64841: outdata = 32'd695;
			64842: outdata = 32'd694;
			64843: outdata = 32'd693;
			64844: outdata = 32'd692;
			64845: outdata = 32'd691;
			64846: outdata = 32'd690;
			64847: outdata = 32'd689;
			64848: outdata = 32'd688;
			64849: outdata = 32'd687;
			64850: outdata = 32'd686;
			64851: outdata = 32'd685;
			64852: outdata = 32'd684;
			64853: outdata = 32'd683;
			64854: outdata = 32'd682;
			64855: outdata = 32'd681;
			64856: outdata = 32'd680;
			64857: outdata = 32'd679;
			64858: outdata = 32'd678;
			64859: outdata = 32'd677;
			64860: outdata = 32'd676;
			64861: outdata = 32'd675;
			64862: outdata = 32'd674;
			64863: outdata = 32'd673;
			64864: outdata = 32'd672;
			64865: outdata = 32'd671;
			64866: outdata = 32'd670;
			64867: outdata = 32'd669;
			64868: outdata = 32'd668;
			64869: outdata = 32'd667;
			64870: outdata = 32'd666;
			64871: outdata = 32'd665;
			64872: outdata = 32'd664;
			64873: outdata = 32'd663;
			64874: outdata = 32'd662;
			64875: outdata = 32'd661;
			64876: outdata = 32'd660;
			64877: outdata = 32'd659;
			64878: outdata = 32'd658;
			64879: outdata = 32'd657;
			64880: outdata = 32'd656;
			64881: outdata = 32'd655;
			64882: outdata = 32'd654;
			64883: outdata = 32'd653;
			64884: outdata = 32'd652;
			64885: outdata = 32'd651;
			64886: outdata = 32'd650;
			64887: outdata = 32'd649;
			64888: outdata = 32'd648;
			64889: outdata = 32'd647;
			64890: outdata = 32'd646;
			64891: outdata = 32'd645;
			64892: outdata = 32'd644;
			64893: outdata = 32'd643;
			64894: outdata = 32'd642;
			64895: outdata = 32'd641;
			64896: outdata = 32'd640;
			64897: outdata = 32'd639;
			64898: outdata = 32'd638;
			64899: outdata = 32'd637;
			64900: outdata = 32'd636;
			64901: outdata = 32'd635;
			64902: outdata = 32'd634;
			64903: outdata = 32'd633;
			64904: outdata = 32'd632;
			64905: outdata = 32'd631;
			64906: outdata = 32'd630;
			64907: outdata = 32'd629;
			64908: outdata = 32'd628;
			64909: outdata = 32'd627;
			64910: outdata = 32'd626;
			64911: outdata = 32'd625;
			64912: outdata = 32'd624;
			64913: outdata = 32'd623;
			64914: outdata = 32'd622;
			64915: outdata = 32'd621;
			64916: outdata = 32'd620;
			64917: outdata = 32'd619;
			64918: outdata = 32'd618;
			64919: outdata = 32'd617;
			64920: outdata = 32'd616;
			64921: outdata = 32'd615;
			64922: outdata = 32'd614;
			64923: outdata = 32'd613;
			64924: outdata = 32'd612;
			64925: outdata = 32'd611;
			64926: outdata = 32'd610;
			64927: outdata = 32'd609;
			64928: outdata = 32'd608;
			64929: outdata = 32'd607;
			64930: outdata = 32'd606;
			64931: outdata = 32'd605;
			64932: outdata = 32'd604;
			64933: outdata = 32'd603;
			64934: outdata = 32'd602;
			64935: outdata = 32'd601;
			64936: outdata = 32'd600;
			64937: outdata = 32'd599;
			64938: outdata = 32'd598;
			64939: outdata = 32'd597;
			64940: outdata = 32'd596;
			64941: outdata = 32'd595;
			64942: outdata = 32'd594;
			64943: outdata = 32'd593;
			64944: outdata = 32'd592;
			64945: outdata = 32'd591;
			64946: outdata = 32'd590;
			64947: outdata = 32'd589;
			64948: outdata = 32'd588;
			64949: outdata = 32'd587;
			64950: outdata = 32'd586;
			64951: outdata = 32'd585;
			64952: outdata = 32'd584;
			64953: outdata = 32'd583;
			64954: outdata = 32'd582;
			64955: outdata = 32'd581;
			64956: outdata = 32'd580;
			64957: outdata = 32'd579;
			64958: outdata = 32'd578;
			64959: outdata = 32'd577;
			64960: outdata = 32'd576;
			64961: outdata = 32'd575;
			64962: outdata = 32'd574;
			64963: outdata = 32'd573;
			64964: outdata = 32'd572;
			64965: outdata = 32'd571;
			64966: outdata = 32'd570;
			64967: outdata = 32'd569;
			64968: outdata = 32'd568;
			64969: outdata = 32'd567;
			64970: outdata = 32'd566;
			64971: outdata = 32'd565;
			64972: outdata = 32'd564;
			64973: outdata = 32'd563;
			64974: outdata = 32'd562;
			64975: outdata = 32'd561;
			64976: outdata = 32'd560;
			64977: outdata = 32'd559;
			64978: outdata = 32'd558;
			64979: outdata = 32'd557;
			64980: outdata = 32'd556;
			64981: outdata = 32'd555;
			64982: outdata = 32'd554;
			64983: outdata = 32'd553;
			64984: outdata = 32'd552;
			64985: outdata = 32'd551;
			64986: outdata = 32'd550;
			64987: outdata = 32'd549;
			64988: outdata = 32'd548;
			64989: outdata = 32'd547;
			64990: outdata = 32'd546;
			64991: outdata = 32'd545;
			64992: outdata = 32'd544;
			64993: outdata = 32'd543;
			64994: outdata = 32'd542;
			64995: outdata = 32'd541;
			64996: outdata = 32'd540;
			64997: outdata = 32'd539;
			64998: outdata = 32'd538;
			64999: outdata = 32'd537;
			65000: outdata = 32'd536;
			65001: outdata = 32'd535;
			65002: outdata = 32'd534;
			65003: outdata = 32'd533;
			65004: outdata = 32'd532;
			65005: outdata = 32'd531;
			65006: outdata = 32'd530;
			65007: outdata = 32'd529;
			65008: outdata = 32'd528;
			65009: outdata = 32'd527;
			65010: outdata = 32'd526;
			65011: outdata = 32'd525;
			65012: outdata = 32'd524;
			65013: outdata = 32'd523;
			65014: outdata = 32'd522;
			65015: outdata = 32'd521;
			65016: outdata = 32'd520;
			65017: outdata = 32'd519;
			65018: outdata = 32'd518;
			65019: outdata = 32'd517;
			65020: outdata = 32'd516;
			65021: outdata = 32'd515;
			65022: outdata = 32'd514;
			65023: outdata = 32'd513;
			65024: outdata = 32'd512;
			65025: outdata = 32'd511;
			65026: outdata = 32'd510;
			65027: outdata = 32'd509;
			65028: outdata = 32'd508;
			65029: outdata = 32'd507;
			65030: outdata = 32'd506;
			65031: outdata = 32'd505;
			65032: outdata = 32'd504;
			65033: outdata = 32'd503;
			65034: outdata = 32'd502;
			65035: outdata = 32'd501;
			65036: outdata = 32'd500;
			65037: outdata = 32'd499;
			65038: outdata = 32'd498;
			65039: outdata = 32'd497;
			65040: outdata = 32'd496;
			65041: outdata = 32'd495;
			65042: outdata = 32'd494;
			65043: outdata = 32'd493;
			65044: outdata = 32'd492;
			65045: outdata = 32'd491;
			65046: outdata = 32'd490;
			65047: outdata = 32'd489;
			65048: outdata = 32'd488;
			65049: outdata = 32'd487;
			65050: outdata = 32'd486;
			65051: outdata = 32'd485;
			65052: outdata = 32'd484;
			65053: outdata = 32'd483;
			65054: outdata = 32'd482;
			65055: outdata = 32'd481;
			65056: outdata = 32'd480;
			65057: outdata = 32'd479;
			65058: outdata = 32'd478;
			65059: outdata = 32'd477;
			65060: outdata = 32'd476;
			65061: outdata = 32'd475;
			65062: outdata = 32'd474;
			65063: outdata = 32'd473;
			65064: outdata = 32'd472;
			65065: outdata = 32'd471;
			65066: outdata = 32'd470;
			65067: outdata = 32'd469;
			65068: outdata = 32'd468;
			65069: outdata = 32'd467;
			65070: outdata = 32'd466;
			65071: outdata = 32'd465;
			65072: outdata = 32'd464;
			65073: outdata = 32'd463;
			65074: outdata = 32'd462;
			65075: outdata = 32'd461;
			65076: outdata = 32'd460;
			65077: outdata = 32'd459;
			65078: outdata = 32'd458;
			65079: outdata = 32'd457;
			65080: outdata = 32'd456;
			65081: outdata = 32'd455;
			65082: outdata = 32'd454;
			65083: outdata = 32'd453;
			65084: outdata = 32'd452;
			65085: outdata = 32'd451;
			65086: outdata = 32'd450;
			65087: outdata = 32'd449;
			65088: outdata = 32'd448;
			65089: outdata = 32'd447;
			65090: outdata = 32'd446;
			65091: outdata = 32'd445;
			65092: outdata = 32'd444;
			65093: outdata = 32'd443;
			65094: outdata = 32'd442;
			65095: outdata = 32'd441;
			65096: outdata = 32'd440;
			65097: outdata = 32'd439;
			65098: outdata = 32'd438;
			65099: outdata = 32'd437;
			65100: outdata = 32'd436;
			65101: outdata = 32'd435;
			65102: outdata = 32'd434;
			65103: outdata = 32'd433;
			65104: outdata = 32'd432;
			65105: outdata = 32'd431;
			65106: outdata = 32'd430;
			65107: outdata = 32'd429;
			65108: outdata = 32'd428;
			65109: outdata = 32'd427;
			65110: outdata = 32'd426;
			65111: outdata = 32'd425;
			65112: outdata = 32'd424;
			65113: outdata = 32'd423;
			65114: outdata = 32'd422;
			65115: outdata = 32'd421;
			65116: outdata = 32'd420;
			65117: outdata = 32'd419;
			65118: outdata = 32'd418;
			65119: outdata = 32'd417;
			65120: outdata = 32'd416;
			65121: outdata = 32'd415;
			65122: outdata = 32'd414;
			65123: outdata = 32'd413;
			65124: outdata = 32'd412;
			65125: outdata = 32'd411;
			65126: outdata = 32'd410;
			65127: outdata = 32'd409;
			65128: outdata = 32'd408;
			65129: outdata = 32'd407;
			65130: outdata = 32'd406;
			65131: outdata = 32'd405;
			65132: outdata = 32'd404;
			65133: outdata = 32'd403;
			65134: outdata = 32'd402;
			65135: outdata = 32'd401;
			65136: outdata = 32'd400;
			65137: outdata = 32'd399;
			65138: outdata = 32'd398;
			65139: outdata = 32'd397;
			65140: outdata = 32'd396;
			65141: outdata = 32'd395;
			65142: outdata = 32'd394;
			65143: outdata = 32'd393;
			65144: outdata = 32'd392;
			65145: outdata = 32'd391;
			65146: outdata = 32'd390;
			65147: outdata = 32'd389;
			65148: outdata = 32'd388;
			65149: outdata = 32'd387;
			65150: outdata = 32'd386;
			65151: outdata = 32'd385;
			65152: outdata = 32'd384;
			65153: outdata = 32'd383;
			65154: outdata = 32'd382;
			65155: outdata = 32'd381;
			65156: outdata = 32'd380;
			65157: outdata = 32'd379;
			65158: outdata = 32'd378;
			65159: outdata = 32'd377;
			65160: outdata = 32'd376;
			65161: outdata = 32'd375;
			65162: outdata = 32'd374;
			65163: outdata = 32'd373;
			65164: outdata = 32'd372;
			65165: outdata = 32'd371;
			65166: outdata = 32'd370;
			65167: outdata = 32'd369;
			65168: outdata = 32'd368;
			65169: outdata = 32'd367;
			65170: outdata = 32'd366;
			65171: outdata = 32'd365;
			65172: outdata = 32'd364;
			65173: outdata = 32'd363;
			65174: outdata = 32'd362;
			65175: outdata = 32'd361;
			65176: outdata = 32'd360;
			65177: outdata = 32'd359;
			65178: outdata = 32'd358;
			65179: outdata = 32'd357;
			65180: outdata = 32'd356;
			65181: outdata = 32'd355;
			65182: outdata = 32'd354;
			65183: outdata = 32'd353;
			65184: outdata = 32'd352;
			65185: outdata = 32'd351;
			65186: outdata = 32'd350;
			65187: outdata = 32'd349;
			65188: outdata = 32'd348;
			65189: outdata = 32'd347;
			65190: outdata = 32'd346;
			65191: outdata = 32'd345;
			65192: outdata = 32'd344;
			65193: outdata = 32'd343;
			65194: outdata = 32'd342;
			65195: outdata = 32'd341;
			65196: outdata = 32'd340;
			65197: outdata = 32'd339;
			65198: outdata = 32'd338;
			65199: outdata = 32'd337;
			65200: outdata = 32'd336;
			65201: outdata = 32'd335;
			65202: outdata = 32'd334;
			65203: outdata = 32'd333;
			65204: outdata = 32'd332;
			65205: outdata = 32'd331;
			65206: outdata = 32'd330;
			65207: outdata = 32'd329;
			65208: outdata = 32'd328;
			65209: outdata = 32'd327;
			65210: outdata = 32'd326;
			65211: outdata = 32'd325;
			65212: outdata = 32'd324;
			65213: outdata = 32'd323;
			65214: outdata = 32'd322;
			65215: outdata = 32'd321;
			65216: outdata = 32'd320;
			65217: outdata = 32'd319;
			65218: outdata = 32'd318;
			65219: outdata = 32'd317;
			65220: outdata = 32'd316;
			65221: outdata = 32'd315;
			65222: outdata = 32'd314;
			65223: outdata = 32'd313;
			65224: outdata = 32'd312;
			65225: outdata = 32'd311;
			65226: outdata = 32'd310;
			65227: outdata = 32'd309;
			65228: outdata = 32'd308;
			65229: outdata = 32'd307;
			65230: outdata = 32'd306;
			65231: outdata = 32'd305;
			65232: outdata = 32'd304;
			65233: outdata = 32'd303;
			65234: outdata = 32'd302;
			65235: outdata = 32'd301;
			65236: outdata = 32'd300;
			65237: outdata = 32'd299;
			65238: outdata = 32'd298;
			65239: outdata = 32'd297;
			65240: outdata = 32'd296;
			65241: outdata = 32'd295;
			65242: outdata = 32'd294;
			65243: outdata = 32'd293;
			65244: outdata = 32'd292;
			65245: outdata = 32'd291;
			65246: outdata = 32'd290;
			65247: outdata = 32'd289;
			65248: outdata = 32'd288;
			65249: outdata = 32'd287;
			65250: outdata = 32'd286;
			65251: outdata = 32'd285;
			65252: outdata = 32'd284;
			65253: outdata = 32'd283;
			65254: outdata = 32'd282;
			65255: outdata = 32'd281;
			65256: outdata = 32'd280;
			65257: outdata = 32'd279;
			65258: outdata = 32'd278;
			65259: outdata = 32'd277;
			65260: outdata = 32'd276;
			65261: outdata = 32'd275;
			65262: outdata = 32'd274;
			65263: outdata = 32'd273;
			65264: outdata = 32'd272;
			65265: outdata = 32'd271;
			65266: outdata = 32'd270;
			65267: outdata = 32'd269;
			65268: outdata = 32'd268;
			65269: outdata = 32'd267;
			65270: outdata = 32'd266;
			65271: outdata = 32'd265;
			65272: outdata = 32'd264;
			65273: outdata = 32'd263;
			65274: outdata = 32'd262;
			65275: outdata = 32'd261;
			65276: outdata = 32'd260;
			65277: outdata = 32'd259;
			65278: outdata = 32'd258;
			65279: outdata = 32'd257;
			65280: outdata = 32'd256;
			65281: outdata = 32'd255;
			65282: outdata = 32'd254;
			65283: outdata = 32'd253;
			65284: outdata = 32'd252;
			65285: outdata = 32'd251;
			65286: outdata = 32'd250;
			65287: outdata = 32'd249;
			65288: outdata = 32'd248;
			65289: outdata = 32'd247;
			65290: outdata = 32'd246;
			65291: outdata = 32'd245;
			65292: outdata = 32'd244;
			65293: outdata = 32'd243;
			65294: outdata = 32'd242;
			65295: outdata = 32'd241;
			65296: outdata = 32'd240;
			65297: outdata = 32'd239;
			65298: outdata = 32'd238;
			65299: outdata = 32'd237;
			65300: outdata = 32'd236;
			65301: outdata = 32'd235;
			65302: outdata = 32'd234;
			65303: outdata = 32'd233;
			65304: outdata = 32'd232;
			65305: outdata = 32'd231;
			65306: outdata = 32'd230;
			65307: outdata = 32'd229;
			65308: outdata = 32'd228;
			65309: outdata = 32'd227;
			65310: outdata = 32'd226;
			65311: outdata = 32'd225;
			65312: outdata = 32'd224;
			65313: outdata = 32'd223;
			65314: outdata = 32'd222;
			65315: outdata = 32'd221;
			65316: outdata = 32'd220;
			65317: outdata = 32'd219;
			65318: outdata = 32'd218;
			65319: outdata = 32'd217;
			65320: outdata = 32'd216;
			65321: outdata = 32'd215;
			65322: outdata = 32'd214;
			65323: outdata = 32'd213;
			65324: outdata = 32'd212;
			65325: outdata = 32'd211;
			65326: outdata = 32'd210;
			65327: outdata = 32'd209;
			65328: outdata = 32'd208;
			65329: outdata = 32'd207;
			65330: outdata = 32'd206;
			65331: outdata = 32'd205;
			65332: outdata = 32'd204;
			65333: outdata = 32'd203;
			65334: outdata = 32'd202;
			65335: outdata = 32'd201;
			65336: outdata = 32'd200;
			65337: outdata = 32'd199;
			65338: outdata = 32'd198;
			65339: outdata = 32'd197;
			65340: outdata = 32'd196;
			65341: outdata = 32'd195;
			65342: outdata = 32'd194;
			65343: outdata = 32'd193;
			65344: outdata = 32'd192;
			65345: outdata = 32'd191;
			65346: outdata = 32'd190;
			65347: outdata = 32'd189;
			65348: outdata = 32'd188;
			65349: outdata = 32'd187;
			65350: outdata = 32'd186;
			65351: outdata = 32'd185;
			65352: outdata = 32'd184;
			65353: outdata = 32'd183;
			65354: outdata = 32'd182;
			65355: outdata = 32'd181;
			65356: outdata = 32'd180;
			65357: outdata = 32'd179;
			65358: outdata = 32'd178;
			65359: outdata = 32'd177;
			65360: outdata = 32'd176;
			65361: outdata = 32'd175;
			65362: outdata = 32'd174;
			65363: outdata = 32'd173;
			65364: outdata = 32'd172;
			65365: outdata = 32'd171;
			65366: outdata = 32'd170;
			65367: outdata = 32'd169;
			65368: outdata = 32'd168;
			65369: outdata = 32'd167;
			65370: outdata = 32'd166;
			65371: outdata = 32'd165;
			65372: outdata = 32'd164;
			65373: outdata = 32'd163;
			65374: outdata = 32'd162;
			65375: outdata = 32'd161;
			65376: outdata = 32'd160;
			65377: outdata = 32'd159;
			65378: outdata = 32'd158;
			65379: outdata = 32'd157;
			65380: outdata = 32'd156;
			65381: outdata = 32'd155;
			65382: outdata = 32'd154;
			65383: outdata = 32'd153;
			65384: outdata = 32'd152;
			65385: outdata = 32'd151;
			65386: outdata = 32'd150;
			65387: outdata = 32'd149;
			65388: outdata = 32'd148;
			65389: outdata = 32'd147;
			65390: outdata = 32'd146;
			65391: outdata = 32'd145;
			65392: outdata = 32'd144;
			65393: outdata = 32'd143;
			65394: outdata = 32'd142;
			65395: outdata = 32'd141;
			65396: outdata = 32'd140;
			65397: outdata = 32'd139;
			65398: outdata = 32'd138;
			65399: outdata = 32'd137;
			65400: outdata = 32'd136;
			65401: outdata = 32'd135;
			65402: outdata = 32'd134;
			65403: outdata = 32'd133;
			65404: outdata = 32'd132;
			65405: outdata = 32'd131;
			65406: outdata = 32'd130;
			65407: outdata = 32'd129;
			65408: outdata = 32'd128;
			65409: outdata = 32'd127;
			65410: outdata = 32'd126;
			65411: outdata = 32'd125;
			65412: outdata = 32'd124;
			65413: outdata = 32'd123;
			65414: outdata = 32'd122;
			65415: outdata = 32'd121;
			65416: outdata = 32'd120;
			65417: outdata = 32'd119;
			65418: outdata = 32'd118;
			65419: outdata = 32'd117;
			65420: outdata = 32'd116;
			65421: outdata = 32'd115;
			65422: outdata = 32'd114;
			65423: outdata = 32'd113;
			65424: outdata = 32'd112;
			65425: outdata = 32'd111;
			65426: outdata = 32'd110;
			65427: outdata = 32'd109;
			65428: outdata = 32'd108;
			65429: outdata = 32'd107;
			65430: outdata = 32'd106;
			65431: outdata = 32'd105;
			65432: outdata = 32'd104;
			65433: outdata = 32'd103;
			65434: outdata = 32'd102;
			65435: outdata = 32'd101;
			65436: outdata = 32'd100;
			65437: outdata = 32'd99;
			65438: outdata = 32'd98;
			65439: outdata = 32'd97;
			65440: outdata = 32'd96;
			65441: outdata = 32'd95;
			65442: outdata = 32'd94;
			65443: outdata = 32'd93;
			65444: outdata = 32'd92;
			65445: outdata = 32'd91;
			65446: outdata = 32'd90;
			65447: outdata = 32'd89;
			65448: outdata = 32'd88;
			65449: outdata = 32'd87;
			65450: outdata = 32'd86;
			65451: outdata = 32'd85;
			65452: outdata = 32'd84;
			65453: outdata = 32'd83;
			65454: outdata = 32'd82;
			65455: outdata = 32'd81;
			65456: outdata = 32'd80;
			65457: outdata = 32'd79;
			65458: outdata = 32'd78;
			65459: outdata = 32'd77;
			65460: outdata = 32'd76;
			65461: outdata = 32'd75;
			65462: outdata = 32'd74;
			65463: outdata = 32'd73;
			65464: outdata = 32'd72;
			65465: outdata = 32'd71;
			65466: outdata = 32'd70;
			65467: outdata = 32'd69;
			65468: outdata = 32'd68;
			65469: outdata = 32'd67;
			65470: outdata = 32'd66;
			65471: outdata = 32'd65;
			65472: outdata = 32'd64;
			65473: outdata = 32'd63;
			65474: outdata = 32'd62;
			65475: outdata = 32'd61;
			65476: outdata = 32'd60;
			65477: outdata = 32'd59;
			65478: outdata = 32'd58;
			65479: outdata = 32'd57;
			65480: outdata = 32'd56;
			65481: outdata = 32'd55;
			65482: outdata = 32'd54;
			65483: outdata = 32'd53;
			65484: outdata = 32'd52;
			65485: outdata = 32'd51;
			65486: outdata = 32'd50;
			65487: outdata = 32'd49;
			65488: outdata = 32'd48;
			65489: outdata = 32'd47;
			65490: outdata = 32'd46;
			65491: outdata = 32'd45;
			65492: outdata = 32'd44;
			65493: outdata = 32'd43;
			65494: outdata = 32'd42;
			65495: outdata = 32'd41;
			65496: outdata = 32'd40;
			65497: outdata = 32'd39;
			65498: outdata = 32'd38;
			65499: outdata = 32'd37;
			65500: outdata = 32'd36;
			65501: outdata = 32'd35;
			65502: outdata = 32'd34;
			65503: outdata = 32'd33;
			65504: outdata = 32'd32;
			65505: outdata = 32'd31;
			65506: outdata = 32'd30;
			65507: outdata = 32'd29;
			65508: outdata = 32'd28;
			65509: outdata = 32'd27;
			65510: outdata = 32'd26;
			65511: outdata = 32'd25;
			65512: outdata = 32'd24;
			65513: outdata = 32'd23;
			65514: outdata = 32'd22;
			65515: outdata = 32'd21;
			65516: outdata = 32'd20;
			65517: outdata = 32'd19;
			65518: outdata = 32'd18;
			65519: outdata = 32'd17;
			65520: outdata = 32'd16;
			65521: outdata = 32'd15;
			65522: outdata = 32'd14;
			65523: outdata = 32'd13;
			65524: outdata = 32'd12;
			65525: outdata = 32'd11;
			65526: outdata = 32'd10;
			65527: outdata = 32'd9;
			65528: outdata = 32'd8;
			65529: outdata = 32'd7;
			65530: outdata = 32'd6;
			65531: outdata = 32'd5;
			65532: outdata = 32'd4;
			65533: outdata = 32'd3;
			65534: outdata = 32'd2;
			65535: outdata = 32'd1;
			default: outdata = 32'b0;
		endcase
	end
endmodule
