module RAM( input [8-1:0] addr, output wire [7:0] outdata );
reg[2039:0] memReg;
	always@(*) begin
		case( addr )
			0: outdata <= memReg[7:0];
			2: outdata <= memReg[15:8];
			3: outdata <= memReg[23:16];
			4: outdata <= memReg[31:24];
			5: outdata <= memReg[39:32];
			6: outdata <= memReg[47:40];
			7: outdata <= memReg[55:48];
			8: outdata <= memReg[63:56];
			9: outdata <= memReg[71:64];
			10: outdata <= memReg[79:72];
			11: outdata <= memReg[87:80];
			12: outdata <= memReg[95:88];
			13: outdata <= memReg[103:96];
			14: outdata <= memReg[111:104];
			15: outdata <= memReg[119:112];
			16: outdata <= memReg[127:120];
			17: outdata <= memReg[135:128];
			18: outdata <= memReg[143:136];
			19: outdata <= memReg[151:144];
			20: outdata <= memReg[159:152];
			21: outdata <= memReg[167:160];
			22: outdata <= memReg[175:168];
			23: outdata <= memReg[183:176];
			24: outdata <= memReg[191:184];
			25: outdata <= memReg[199:192];
			26: outdata <= memReg[207:200];
			27: outdata <= memReg[215:208];
			28: outdata <= memReg[223:216];
			29: outdata <= memReg[231:224];
			30: outdata <= memReg[239:232];
			31: outdata <= memReg[247:240];
			32: outdata <= memReg[255:248];
			33: outdata <= memReg[263:256];
			34: outdata <= memReg[271:264];
			35: outdata <= memReg[279:272];
			36: outdata <= memReg[287:280];
			37: outdata <= memReg[295:288];
			38: outdata <= memReg[303:296];
			39: outdata <= memReg[311:304];
			40: outdata <= memReg[319:312];
			41: outdata <= memReg[327:320];
			42: outdata <= memReg[335:328];
			43: outdata <= memReg[343:336];
			44: outdata <= memReg[351:344];
			45: outdata <= memReg[359:352];
			46: outdata <= memReg[367:360];
			47: outdata <= memReg[375:368];
			48: outdata <= memReg[383:376];
			49: outdata <= memReg[391:384];
			50: outdata <= memReg[399:392];
			51: outdata <= memReg[407:400];
			52: outdata <= memReg[415:408];
			53: outdata <= memReg[423:416];
			54: outdata <= memReg[431:424];
			55: outdata <= memReg[439:432];
			56: outdata <= memReg[447:440];
			57: outdata <= memReg[455:448];
			58: outdata <= memReg[463:456];
			59: outdata <= memReg[471:464];
			60: outdata <= memReg[479:472];
			61: outdata <= memReg[487:480];
			62: outdata <= memReg[495:488];
			63: outdata <= memReg[503:496];
			64: outdata <= memReg[511:504];
			65: outdata <= memReg[519:512];
			66: outdata <= memReg[527:520];
			67: outdata <= memReg[535:528];
			68: outdata <= memReg[543:536];
			69: outdata <= memReg[551:544];
			70: outdata <= memReg[559:552];
			71: outdata <= memReg[567:560];
			72: outdata <= memReg[575:568];
			73: outdata <= memReg[583:576];
			74: outdata <= memReg[591:584];
			75: outdata <= memReg[599:592];
			76: outdata <= memReg[607:600];
			77: outdata <= memReg[615:608];
			78: outdata <= memReg[623:616];
			79: outdata <= memReg[631:624];
			80: outdata <= memReg[639:632];
			81: outdata <= memReg[647:640];
			82: outdata <= memReg[655:648];
			83: outdata <= memReg[663:656];
			84: outdata <= memReg[671:664];
			85: outdata <= memReg[679:672];
			86: outdata <= memReg[687:680];
			87: outdata <= memReg[695:688];
			88: outdata <= memReg[703:696];
			89: outdata <= memReg[711:704];
			90: outdata <= memReg[719:712];
			91: outdata <= memReg[727:720];
			92: outdata <= memReg[735:728];
			93: outdata <= memReg[743:736];
			94: outdata <= memReg[751:744];
			95: outdata <= memReg[759:752];
			96: outdata <= memReg[767:760];
			97: outdata <= memReg[775:768];
			98: outdata <= memReg[783:776];
			99: outdata <= memReg[791:784];
			100: outdata <= memReg[799:792];
			101: outdata <= memReg[807:800];
			102: outdata <= memReg[815:808];
			103: outdata <= memReg[823:816];
			104: outdata <= memReg[831:824];
			105: outdata <= memReg[839:832];
			106: outdata <= memReg[847:840];
			107: outdata <= memReg[855:848];
			108: outdata <= memReg[863:856];
			109: outdata <= memReg[871:864];
			110: outdata <= memReg[879:872];
			111: outdata <= memReg[887:880];
			112: outdata <= memReg[895:888];
			113: outdata <= memReg[903:896];
			114: outdata <= memReg[911:904];
			115: outdata <= memReg[919:912];
			116: outdata <= memReg[927:920];
			117: outdata <= memReg[935:928];
			118: outdata <= memReg[943:936];
			119: outdata <= memReg[951:944];
			120: outdata <= memReg[959:952];
			121: outdata <= memReg[967:960];
			122: outdata <= memReg[975:968];
			123: outdata <= memReg[983:976];
			124: outdata <= memReg[991:984];
			125: outdata <= memReg[999:992];
			126: outdata <= memReg[1007:1000];
			127: outdata <= memReg[1015:1008];
			128: outdata <= memReg[1023:1016];
			129: outdata <= memReg[1031:1024];
			130: outdata <= memReg[1039:1032];
			131: outdata <= memReg[1047:1040];
			132: outdata <= memReg[1055:1048];
			133: outdata <= memReg[1063:1056];
			134: outdata <= memReg[1071:1064];
			135: outdata <= memReg[1079:1072];
			136: outdata <= memReg[1087:1080];
			137: outdata <= memReg[1095:1088];
			138: outdata <= memReg[1103:1096];
			139: outdata <= memReg[1111:1104];
			140: outdata <= memReg[1119:1112];
			141: outdata <= memReg[1127:1120];
			142: outdata <= memReg[1135:1128];
			143: outdata <= memReg[1143:1136];
			144: outdata <= memReg[1151:1144];
			145: outdata <= memReg[1159:1152];
			146: outdata <= memReg[1167:1160];
			147: outdata <= memReg[1175:1168];
			148: outdata <= memReg[1183:1176];
			149: outdata <= memReg[1191:1184];
			150: outdata <= memReg[1199:1192];
			151: outdata <= memReg[1207:1200];
			152: outdata <= memReg[1215:1208];
			153: outdata <= memReg[1223:1216];
			154: outdata <= memReg[1231:1224];
			155: outdata <= memReg[1239:1232];
			156: outdata <= memReg[1247:1240];
			157: outdata <= memReg[1255:1248];
			158: outdata <= memReg[1263:1256];
			159: outdata <= memReg[1271:1264];
			160: outdata <= memReg[1279:1272];
			161: outdata <= memReg[1287:1280];
			162: outdata <= memReg[1295:1288];
			163: outdata <= memReg[1303:1296];
			164: outdata <= memReg[1311:1304];
			165: outdata <= memReg[1319:1312];
			166: outdata <= memReg[1327:1320];
			167: outdata <= memReg[1335:1328];
			168: outdata <= memReg[1343:1336];
			169: outdata <= memReg[1351:1344];
			170: outdata <= memReg[1359:1352];
			171: outdata <= memReg[1367:1360];
			172: outdata <= memReg[1375:1368];
			173: outdata <= memReg[1383:1376];
			174: outdata <= memReg[1391:1384];
			175: outdata <= memReg[1399:1392];
			176: outdata <= memReg[1407:1400];
			177: outdata <= memReg[1415:1408];
			178: outdata <= memReg[1423:1416];
			179: outdata <= memReg[1431:1424];
			180: outdata <= memReg[1439:1432];
			181: outdata <= memReg[1447:1440];
			182: outdata <= memReg[1455:1448];
			183: outdata <= memReg[1463:1456];
			184: outdata <= memReg[1471:1464];
			185: outdata <= memReg[1479:1472];
			186: outdata <= memReg[1487:1480];
			187: outdata <= memReg[1495:1488];
			188: outdata <= memReg[1503:1496];
			189: outdata <= memReg[1511:1504];
			190: outdata <= memReg[1519:1512];
			191: outdata <= memReg[1527:1520];
			192: outdata <= memReg[1535:1528];
			193: outdata <= memReg[1543:1536];
			194: outdata <= memReg[1551:1544];
			195: outdata <= memReg[1559:1552];
			196: outdata <= memReg[1567:1560];
			197: outdata <= memReg[1575:1568];
			198: outdata <= memReg[1583:1576];
			199: outdata <= memReg[1591:1584];
			200: outdata <= memReg[1599:1592];
			201: outdata <= memReg[1607:1600];
			202: outdata <= memReg[1615:1608];
			203: outdata <= memReg[1623:1616];
			204: outdata <= memReg[1631:1624];
			205: outdata <= memReg[1639:1632];
			206: outdata <= memReg[1647:1640];
			207: outdata <= memReg[1655:1648];
			208: outdata <= memReg[1663:1656];
			209: outdata <= memReg[1671:1664];
			210: outdata <= memReg[1679:1672];
			211: outdata <= memReg[1687:1680];
			212: outdata <= memReg[1695:1688];
			213: outdata <= memReg[1703:1696];
			214: outdata <= memReg[1711:1704];
			215: outdata <= memReg[1719:1712];
			216: outdata <= memReg[1727:1720];
			217: outdata <= memReg[1735:1728];
			218: outdata <= memReg[1743:1736];
			219: outdata <= memReg[1751:1744];
			220: outdata <= memReg[1759:1752];
			221: outdata <= memReg[1767:1760];
			222: outdata <= memReg[1775:1768];
			223: outdata <= memReg[1783:1776];
			224: outdata <= memReg[1791:1784];
			225: outdata <= memReg[1799:1792];
			226: outdata <= memReg[1807:1800];
			227: outdata <= memReg[1815:1808];
			228: outdata <= memReg[1823:1816];
			229: outdata <= memReg[1831:1824];
			230: outdata <= memReg[1839:1832];
			231: outdata <= memReg[1847:1840];
			232: outdata <= memReg[1855:1848];
			233: outdata <= memReg[1863:1856];
			234: outdata <= memReg[1871:1864];
			235: outdata <= memReg[1879:1872];
			236: outdata <= memReg[1887:1880];
			237: outdata <= memReg[1895:1888];
			238: outdata <= memReg[1903:1896];
			239: outdata <= memReg[1911:1904];
			240: outdata <= memReg[1919:1912];
			241: outdata <= memReg[1927:1920];
			242: outdata <= memReg[1935:1928];
			243: outdata <= memReg[1943:1936];
			244: outdata <= memReg[1951:1944];
			245: outdata <= memReg[1959:1952];
			246: outdata <= memReg[1967:1960];
			247: outdata <= memReg[1975:1968];
			248: outdata <= memReg[1983:1976];
			249: outdata <= memReg[1991:1984];
			250: outdata <= memReg[1999:1992];
			251: outdata <= memReg[2007:2000];
			252: outdata <= memReg[2015:2008];
			253: outdata <= memReg[2023:2016];
			254: outdata <= memReg[2031:2024];
			255: outdata <= memReg[2039:2032];
			default: outdata <= 8'b0;
		endcase
	end
endmodule
